VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO TopModule
  CLASS BLOCK ;
  FOREIGN TopModule ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 28.940 10.640 30.540 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 182.540 10.640 184.140 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 336.140 10.640 337.740 389.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 30.030 389.860 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 183.210 389.860 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 336.390 389.860 337.990 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 25.640 10.640 27.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 179.240 10.640 180.840 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.840 10.640 334.440 389.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 26.730 389.860 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 179.910 389.860 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 9.880 333.090 389.860 334.690 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END clk
  PIN ctrl[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END ctrl[0]
  PIN ctrl[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END ctrl[1]
  PIN data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.840 400.000 194.440 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 396.000 293.390 400.000 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 258.440 400.000 259.040 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 187.040 400.000 187.640 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 396.000 119.510 400.000 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 396.000 200.010 400.000 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 396.000 270.850 400.000 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 105.440 400.000 106.040 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 183.640 400.000 184.240 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 396.000 209.670 400.000 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 396.000 190.440 400.000 191.040 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 396.000 248.310 400.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 248.240 400.000 248.840 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 396.000 164.590 400.000 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 81.640 400.000 82.240 ;
    END
  END data_out[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.040 400.000 170.640 ;
    END
  END reset
  OBS
      LAYER nwell ;
        RECT 9.930 10.795 389.810 389.150 ;
      LAYER li1 ;
        RECT 10.120 10.795 389.620 389.045 ;
      LAYER met1 ;
        RECT 6.050 10.640 389.620 389.200 ;
      LAYER met2 ;
        RECT 6.070 395.720 118.950 396.000 ;
        RECT 119.790 395.720 164.030 396.000 ;
        RECT 164.870 395.720 199.450 396.000 ;
        RECT 200.290 395.720 209.110 396.000 ;
        RECT 209.950 395.720 247.750 396.000 ;
        RECT 248.590 395.720 270.290 396.000 ;
        RECT 271.130 395.720 292.830 396.000 ;
        RECT 293.670 395.720 388.150 396.000 ;
        RECT 6.070 4.280 388.150 395.720 ;
        RECT 6.070 4.000 112.510 4.280 ;
        RECT 113.350 4.000 115.730 4.280 ;
        RECT 116.570 4.000 167.250 4.280 ;
        RECT 168.090 4.000 209.110 4.280 ;
        RECT 209.950 4.000 212.330 4.280 ;
        RECT 213.170 4.000 221.990 4.280 ;
        RECT 222.830 4.000 260.630 4.280 ;
        RECT 261.470 4.000 289.610 4.280 ;
        RECT 290.450 4.000 296.050 4.280 ;
        RECT 296.890 4.000 388.150 4.280 ;
      LAYER met3 ;
        RECT 4.000 259.440 396.000 389.125 ;
        RECT 4.000 258.040 395.600 259.440 ;
        RECT 4.000 249.240 396.000 258.040 ;
        RECT 4.000 247.840 395.600 249.240 ;
        RECT 4.000 228.840 396.000 247.840 ;
        RECT 4.400 227.440 396.000 228.840 ;
        RECT 4.000 208.440 396.000 227.440 ;
        RECT 4.400 207.040 396.000 208.440 ;
        RECT 4.000 194.840 396.000 207.040 ;
        RECT 4.000 193.440 395.600 194.840 ;
        RECT 4.000 191.440 396.000 193.440 ;
        RECT 4.000 190.040 395.600 191.440 ;
        RECT 4.000 188.040 396.000 190.040 ;
        RECT 4.000 186.640 395.600 188.040 ;
        RECT 4.000 184.640 396.000 186.640 ;
        RECT 4.000 183.240 395.600 184.640 ;
        RECT 4.000 177.840 396.000 183.240 ;
        RECT 4.400 176.440 396.000 177.840 ;
        RECT 4.000 171.040 396.000 176.440 ;
        RECT 4.000 169.640 395.600 171.040 ;
        RECT 4.000 160.840 396.000 169.640 ;
        RECT 4.400 159.440 396.000 160.840 ;
        RECT 4.000 143.840 396.000 159.440 ;
        RECT 4.400 142.440 396.000 143.840 ;
        RECT 4.000 140.440 396.000 142.440 ;
        RECT 4.400 139.040 396.000 140.440 ;
        RECT 4.000 133.640 396.000 139.040 ;
        RECT 4.400 132.240 396.000 133.640 ;
        RECT 4.000 130.240 396.000 132.240 ;
        RECT 4.400 128.840 396.000 130.240 ;
        RECT 4.000 116.640 396.000 128.840 ;
        RECT 4.400 115.240 396.000 116.640 ;
        RECT 4.000 106.440 396.000 115.240 ;
        RECT 4.000 105.040 395.600 106.440 ;
        RECT 4.000 82.640 396.000 105.040 ;
        RECT 4.000 81.240 395.600 82.640 ;
        RECT 4.000 10.715 396.000 81.240 ;
  END
END TopModule
END LIBRARY

