magic
tech sky130A
magscale 1 2
timestamp 1749953730
<< viali >>
rect 23949 77673 23983 77707
rect 33057 77673 33091 77707
rect 40049 77673 40083 77707
rect 41981 77673 42015 77707
rect 49709 77673 49743 77707
rect 54217 77673 54251 77707
rect 58817 77673 58851 77707
rect 77585 51765 77619 51799
rect 77585 49725 77619 49759
rect 64889 43809 64923 43843
rect 64981 43741 65015 43775
rect 66545 43741 66579 43775
rect 67097 43741 67131 43775
rect 65349 43605 65383 43639
rect 66913 43401 66947 43435
rect 65441 43333 65475 43367
rect 67097 43333 67131 43367
rect 67189 43265 67223 43299
rect 65165 43197 65199 43231
rect 59369 42721 59403 42755
rect 60105 42721 60139 42755
rect 57621 42653 57655 42687
rect 57897 42585 57931 42619
rect 59553 42517 59587 42551
rect 58081 42313 58115 42347
rect 58909 42313 58943 42347
rect 58173 42177 58207 42211
rect 59001 42177 59035 42211
rect 64705 41769 64739 41803
rect 2329 41565 2363 41599
rect 64613 41565 64647 41599
rect 64797 41565 64831 41599
rect 71329 41565 71363 41599
rect 74365 41565 74399 41599
rect 76389 41565 76423 41599
rect 74641 41497 74675 41531
rect 76297 41497 76331 41531
rect 71237 41429 71271 41463
rect 76113 41429 76147 41463
rect 70225 41089 70259 41123
rect 74457 41089 74491 41123
rect 75285 41089 75319 41123
rect 70501 41021 70535 41055
rect 74365 41021 74399 41055
rect 74825 41021 74859 41055
rect 75929 41021 75963 41055
rect 71973 40885 72007 40919
rect 61209 40681 61243 40715
rect 61650 40681 61684 40715
rect 70685 40681 70719 40715
rect 63141 40613 63175 40647
rect 66545 40613 66579 40647
rect 70869 40613 70903 40647
rect 60933 40545 60967 40579
rect 65901 40545 65935 40579
rect 68293 40545 68327 40579
rect 71145 40545 71179 40579
rect 60841 40477 60875 40511
rect 61393 40477 61427 40511
rect 65809 40477 65843 40511
rect 65993 40477 66027 40511
rect 66085 40477 66119 40511
rect 68017 40409 68051 40443
rect 66269 40341 66303 40375
rect 62037 40137 62071 40171
rect 65809 40137 65843 40171
rect 66729 40137 66763 40171
rect 65901 40069 65935 40103
rect 66177 40069 66211 40103
rect 61761 40001 61795 40035
rect 61853 40001 61887 40035
rect 62681 40001 62715 40035
rect 65993 40001 66027 40035
rect 67189 40001 67223 40035
rect 67281 40001 67315 40035
rect 66269 39933 66303 39967
rect 66545 39865 66579 39899
rect 65625 39797 65659 39831
rect 70869 39593 70903 39627
rect 66545 39525 66579 39559
rect 76205 39525 76239 39559
rect 56793 39457 56827 39491
rect 58817 39389 58851 39423
rect 66729 39389 66763 39423
rect 66821 39389 66855 39423
rect 75929 39389 75963 39423
rect 57069 39321 57103 39355
rect 58725 39321 58759 39355
rect 71145 39321 71179 39355
rect 71421 39321 71455 39355
rect 76205 39321 76239 39355
rect 58541 39253 58575 39287
rect 66913 39253 66947 39287
rect 67097 39253 67131 39287
rect 71053 39253 71087 39287
rect 71237 39253 71271 39287
rect 76021 39253 76055 39287
rect 71145 39049 71179 39083
rect 71513 39049 71547 39083
rect 71605 39049 71639 39083
rect 75469 39049 75503 39083
rect 65441 38913 65475 38947
rect 70869 38913 70903 38947
rect 71237 38913 71271 38947
rect 71789 38913 71823 38947
rect 71973 38913 72007 38947
rect 75561 38913 75595 38947
rect 77309 38913 77343 38947
rect 70961 38845 70995 38879
rect 71329 38845 71363 38879
rect 75377 38845 75411 38879
rect 77493 38777 77527 38811
rect 66729 38709 66763 38743
rect 75929 38709 75963 38743
rect 57069 38505 57103 38539
rect 63417 38505 63451 38539
rect 69121 38505 69155 38539
rect 74733 38505 74767 38539
rect 76297 38505 76331 38539
rect 57253 38301 57287 38335
rect 57345 38301 57379 38335
rect 74641 38301 74675 38335
rect 76113 38301 76147 38335
rect 77309 38301 77343 38335
rect 57621 38233 57655 38267
rect 57805 38233 57839 38267
rect 57989 38233 58023 38267
rect 64705 38233 64739 38267
rect 67833 38233 67867 38267
rect 77493 38165 77527 38199
rect 67925 37893 67959 37927
rect 77309 37825 77343 37859
rect 77493 37621 77527 37655
rect 64337 37281 64371 37315
rect 64613 37281 64647 37315
rect 57529 37213 57563 37247
rect 57713 37213 57747 37247
rect 67097 37213 67131 37247
rect 75377 37213 75411 37247
rect 77309 37213 77343 37247
rect 75285 37145 75319 37179
rect 57621 37077 57655 37111
rect 66085 37077 66119 37111
rect 66545 37077 66579 37111
rect 77493 37077 77527 37111
rect 65441 36873 65475 36907
rect 66085 36873 66119 36907
rect 60013 36805 60047 36839
rect 60381 36805 60415 36839
rect 60749 36805 60783 36839
rect 60197 36737 60231 36771
rect 60289 36737 60323 36771
rect 65625 36737 65659 36771
rect 65809 36737 65843 36771
rect 65901 36737 65935 36771
rect 66177 36737 66211 36771
rect 66637 36329 66671 36363
rect 76481 36329 76515 36363
rect 60473 36261 60507 36295
rect 60657 36261 60691 36295
rect 70777 36261 70811 36295
rect 60105 36193 60139 36227
rect 60197 36193 60231 36227
rect 60289 36193 60323 36227
rect 61025 36193 61059 36227
rect 72709 36193 72743 36227
rect 60013 36125 60047 36159
rect 66545 36125 66579 36159
rect 66729 36125 66763 36159
rect 70593 36125 70627 36159
rect 70869 36125 70903 36159
rect 72801 36125 72835 36159
rect 74089 36125 74123 36159
rect 76205 36125 76239 36159
rect 76297 36125 76331 36159
rect 70685 36057 70719 36091
rect 74365 36057 74399 36091
rect 76113 36057 76147 36091
rect 60565 35989 60599 36023
rect 73169 35989 73203 36023
rect 75837 35989 75871 36023
rect 74365 35785 74399 35819
rect 60657 35717 60691 35751
rect 62313 35717 62347 35751
rect 56701 35649 56735 35683
rect 57437 35649 57471 35683
rect 58081 35649 58115 35683
rect 62405 35649 62439 35683
rect 71145 35649 71179 35683
rect 71237 35649 71271 35683
rect 71697 35649 71731 35683
rect 75009 35649 75043 35683
rect 56793 35581 56827 35615
rect 60381 35581 60415 35615
rect 62129 35581 62163 35615
rect 70133 35581 70167 35615
rect 70777 35581 70811 35615
rect 70961 35581 70995 35615
rect 71053 35581 71087 35615
rect 71421 35581 71455 35615
rect 71881 35581 71915 35615
rect 2329 35445 2363 35479
rect 56425 35445 56459 35479
rect 71513 35445 71547 35479
rect 56590 35241 56624 35275
rect 58081 35241 58115 35275
rect 70961 35241 70995 35275
rect 56333 35105 56367 35139
rect 58357 35037 58391 35071
rect 70685 35037 70719 35071
rect 70777 35037 70811 35071
rect 58265 34969 58299 35003
rect 71329 34629 71363 34663
rect 77309 34629 77343 34663
rect 65901 34561 65935 34595
rect 66361 34561 66395 34595
rect 67005 34561 67039 34595
rect 71605 34561 71639 34595
rect 72157 34561 72191 34595
rect 77493 34561 77527 34595
rect 65993 34493 66027 34527
rect 69857 34493 69891 34527
rect 71881 34493 71915 34527
rect 66177 34357 66211 34391
rect 66545 34153 66579 34187
rect 70961 34153 70995 34187
rect 68017 34017 68051 34051
rect 68293 34017 68327 34051
rect 71053 33949 71087 33983
rect 66913 33609 66947 33643
rect 66821 33473 66855 33507
rect 2329 32181 2363 32215
rect 2329 28985 2363 29019
rect 2329 27965 2363 27999
rect 2329 26741 2363 26775
rect 2329 26333 2363 26367
rect 2329 23477 2363 23511
rect 77585 21301 77619 21335
rect 77585 16609 77619 16643
rect 22753 2397 22787 2431
rect 23305 2397 23339 2431
rect 33609 2397 33643 2431
rect 41981 2397 42015 2431
rect 42625 2397 42659 2431
rect 44557 2397 44591 2431
rect 52285 2397 52319 2431
rect 58081 2397 58115 2431
rect 59369 2397 59403 2431
<< metal1 >>
rect 2024 77818 77924 77840
rect 2024 77766 5134 77818
rect 5186 77766 5198 77818
rect 5250 77766 5262 77818
rect 5314 77766 5326 77818
rect 5378 77766 5390 77818
rect 5442 77766 35854 77818
rect 35906 77766 35918 77818
rect 35970 77766 35982 77818
rect 36034 77766 36046 77818
rect 36098 77766 36110 77818
rect 36162 77766 66574 77818
rect 66626 77766 66638 77818
rect 66690 77766 66702 77818
rect 66754 77766 66766 77818
rect 66818 77766 66830 77818
rect 66882 77766 77924 77818
rect 2024 77744 77924 77766
rect 23842 77664 23848 77716
rect 23900 77704 23906 77716
rect 23937 77707 23995 77713
rect 23937 77704 23949 77707
rect 23900 77676 23949 77704
rect 23900 77664 23906 77676
rect 23937 77673 23949 77676
rect 23983 77673 23995 77707
rect 23937 77667 23995 77673
rect 32858 77664 32864 77716
rect 32916 77704 32922 77716
rect 33045 77707 33103 77713
rect 33045 77704 33057 77707
rect 32916 77676 33057 77704
rect 32916 77664 32922 77676
rect 33045 77673 33057 77676
rect 33091 77673 33103 77707
rect 33045 77667 33103 77673
rect 39942 77664 39948 77716
rect 40000 77704 40006 77716
rect 40037 77707 40095 77713
rect 40037 77704 40049 77707
rect 40000 77676 40049 77704
rect 40000 77664 40006 77676
rect 40037 77673 40049 77676
rect 40083 77673 40095 77707
rect 40037 77667 40095 77673
rect 41874 77664 41880 77716
rect 41932 77704 41938 77716
rect 41969 77707 42027 77713
rect 41969 77704 41981 77707
rect 41932 77676 41981 77704
rect 41932 77664 41938 77676
rect 41969 77673 41981 77676
rect 42015 77673 42027 77707
rect 41969 77667 42027 77673
rect 49602 77664 49608 77716
rect 49660 77704 49666 77716
rect 49697 77707 49755 77713
rect 49697 77704 49709 77707
rect 49660 77676 49709 77704
rect 49660 77664 49666 77676
rect 49697 77673 49709 77676
rect 49743 77673 49755 77707
rect 49697 77667 49755 77673
rect 54110 77664 54116 77716
rect 54168 77704 54174 77716
rect 54205 77707 54263 77713
rect 54205 77704 54217 77707
rect 54168 77676 54217 77704
rect 54168 77664 54174 77676
rect 54205 77673 54217 77676
rect 54251 77673 54263 77707
rect 54205 77667 54263 77673
rect 58618 77664 58624 77716
rect 58676 77704 58682 77716
rect 58805 77707 58863 77713
rect 58805 77704 58817 77707
rect 58676 77676 58817 77704
rect 58676 77664 58682 77676
rect 58805 77673 58817 77676
rect 58851 77673 58863 77707
rect 58805 77667 58863 77673
rect 2024 77274 77924 77296
rect 2024 77222 5794 77274
rect 5846 77222 5858 77274
rect 5910 77222 5922 77274
rect 5974 77222 5986 77274
rect 6038 77222 6050 77274
rect 6102 77222 36514 77274
rect 36566 77222 36578 77274
rect 36630 77222 36642 77274
rect 36694 77222 36706 77274
rect 36758 77222 36770 77274
rect 36822 77222 67234 77274
rect 67286 77222 67298 77274
rect 67350 77222 67362 77274
rect 67414 77222 67426 77274
rect 67478 77222 67490 77274
rect 67542 77222 77924 77274
rect 2024 77200 77924 77222
rect 2024 76730 77924 76752
rect 2024 76678 5134 76730
rect 5186 76678 5198 76730
rect 5250 76678 5262 76730
rect 5314 76678 5326 76730
rect 5378 76678 5390 76730
rect 5442 76678 35854 76730
rect 35906 76678 35918 76730
rect 35970 76678 35982 76730
rect 36034 76678 36046 76730
rect 36098 76678 36110 76730
rect 36162 76678 66574 76730
rect 66626 76678 66638 76730
rect 66690 76678 66702 76730
rect 66754 76678 66766 76730
rect 66818 76678 66830 76730
rect 66882 76678 77924 76730
rect 2024 76656 77924 76678
rect 2024 76186 77924 76208
rect 2024 76134 5794 76186
rect 5846 76134 5858 76186
rect 5910 76134 5922 76186
rect 5974 76134 5986 76186
rect 6038 76134 6050 76186
rect 6102 76134 36514 76186
rect 36566 76134 36578 76186
rect 36630 76134 36642 76186
rect 36694 76134 36706 76186
rect 36758 76134 36770 76186
rect 36822 76134 67234 76186
rect 67286 76134 67298 76186
rect 67350 76134 67362 76186
rect 67414 76134 67426 76186
rect 67478 76134 67490 76186
rect 67542 76134 77924 76186
rect 2024 76112 77924 76134
rect 2024 75642 77924 75664
rect 2024 75590 5134 75642
rect 5186 75590 5198 75642
rect 5250 75590 5262 75642
rect 5314 75590 5326 75642
rect 5378 75590 5390 75642
rect 5442 75590 35854 75642
rect 35906 75590 35918 75642
rect 35970 75590 35982 75642
rect 36034 75590 36046 75642
rect 36098 75590 36110 75642
rect 36162 75590 66574 75642
rect 66626 75590 66638 75642
rect 66690 75590 66702 75642
rect 66754 75590 66766 75642
rect 66818 75590 66830 75642
rect 66882 75590 77924 75642
rect 2024 75568 77924 75590
rect 2024 75098 77924 75120
rect 2024 75046 5794 75098
rect 5846 75046 5858 75098
rect 5910 75046 5922 75098
rect 5974 75046 5986 75098
rect 6038 75046 6050 75098
rect 6102 75046 36514 75098
rect 36566 75046 36578 75098
rect 36630 75046 36642 75098
rect 36694 75046 36706 75098
rect 36758 75046 36770 75098
rect 36822 75046 67234 75098
rect 67286 75046 67298 75098
rect 67350 75046 67362 75098
rect 67414 75046 67426 75098
rect 67478 75046 67490 75098
rect 67542 75046 77924 75098
rect 2024 75024 77924 75046
rect 2024 74554 77924 74576
rect 2024 74502 5134 74554
rect 5186 74502 5198 74554
rect 5250 74502 5262 74554
rect 5314 74502 5326 74554
rect 5378 74502 5390 74554
rect 5442 74502 35854 74554
rect 35906 74502 35918 74554
rect 35970 74502 35982 74554
rect 36034 74502 36046 74554
rect 36098 74502 36110 74554
rect 36162 74502 66574 74554
rect 66626 74502 66638 74554
rect 66690 74502 66702 74554
rect 66754 74502 66766 74554
rect 66818 74502 66830 74554
rect 66882 74502 77924 74554
rect 2024 74480 77924 74502
rect 2024 74010 77924 74032
rect 2024 73958 5794 74010
rect 5846 73958 5858 74010
rect 5910 73958 5922 74010
rect 5974 73958 5986 74010
rect 6038 73958 6050 74010
rect 6102 73958 36514 74010
rect 36566 73958 36578 74010
rect 36630 73958 36642 74010
rect 36694 73958 36706 74010
rect 36758 73958 36770 74010
rect 36822 73958 67234 74010
rect 67286 73958 67298 74010
rect 67350 73958 67362 74010
rect 67414 73958 67426 74010
rect 67478 73958 67490 74010
rect 67542 73958 77924 74010
rect 2024 73936 77924 73958
rect 2024 73466 77924 73488
rect 2024 73414 5134 73466
rect 5186 73414 5198 73466
rect 5250 73414 5262 73466
rect 5314 73414 5326 73466
rect 5378 73414 5390 73466
rect 5442 73414 35854 73466
rect 35906 73414 35918 73466
rect 35970 73414 35982 73466
rect 36034 73414 36046 73466
rect 36098 73414 36110 73466
rect 36162 73414 66574 73466
rect 66626 73414 66638 73466
rect 66690 73414 66702 73466
rect 66754 73414 66766 73466
rect 66818 73414 66830 73466
rect 66882 73414 77924 73466
rect 2024 73392 77924 73414
rect 2024 72922 77924 72944
rect 2024 72870 5794 72922
rect 5846 72870 5858 72922
rect 5910 72870 5922 72922
rect 5974 72870 5986 72922
rect 6038 72870 6050 72922
rect 6102 72870 36514 72922
rect 36566 72870 36578 72922
rect 36630 72870 36642 72922
rect 36694 72870 36706 72922
rect 36758 72870 36770 72922
rect 36822 72870 67234 72922
rect 67286 72870 67298 72922
rect 67350 72870 67362 72922
rect 67414 72870 67426 72922
rect 67478 72870 67490 72922
rect 67542 72870 77924 72922
rect 2024 72848 77924 72870
rect 2024 72378 77924 72400
rect 2024 72326 5134 72378
rect 5186 72326 5198 72378
rect 5250 72326 5262 72378
rect 5314 72326 5326 72378
rect 5378 72326 5390 72378
rect 5442 72326 35854 72378
rect 35906 72326 35918 72378
rect 35970 72326 35982 72378
rect 36034 72326 36046 72378
rect 36098 72326 36110 72378
rect 36162 72326 66574 72378
rect 66626 72326 66638 72378
rect 66690 72326 66702 72378
rect 66754 72326 66766 72378
rect 66818 72326 66830 72378
rect 66882 72326 77924 72378
rect 2024 72304 77924 72326
rect 2024 71834 77924 71856
rect 2024 71782 5794 71834
rect 5846 71782 5858 71834
rect 5910 71782 5922 71834
rect 5974 71782 5986 71834
rect 6038 71782 6050 71834
rect 6102 71782 36514 71834
rect 36566 71782 36578 71834
rect 36630 71782 36642 71834
rect 36694 71782 36706 71834
rect 36758 71782 36770 71834
rect 36822 71782 67234 71834
rect 67286 71782 67298 71834
rect 67350 71782 67362 71834
rect 67414 71782 67426 71834
rect 67478 71782 67490 71834
rect 67542 71782 77924 71834
rect 2024 71760 77924 71782
rect 2024 71290 77924 71312
rect 2024 71238 5134 71290
rect 5186 71238 5198 71290
rect 5250 71238 5262 71290
rect 5314 71238 5326 71290
rect 5378 71238 5390 71290
rect 5442 71238 35854 71290
rect 35906 71238 35918 71290
rect 35970 71238 35982 71290
rect 36034 71238 36046 71290
rect 36098 71238 36110 71290
rect 36162 71238 66574 71290
rect 66626 71238 66638 71290
rect 66690 71238 66702 71290
rect 66754 71238 66766 71290
rect 66818 71238 66830 71290
rect 66882 71238 77924 71290
rect 2024 71216 77924 71238
rect 2024 70746 77924 70768
rect 2024 70694 5794 70746
rect 5846 70694 5858 70746
rect 5910 70694 5922 70746
rect 5974 70694 5986 70746
rect 6038 70694 6050 70746
rect 6102 70694 36514 70746
rect 36566 70694 36578 70746
rect 36630 70694 36642 70746
rect 36694 70694 36706 70746
rect 36758 70694 36770 70746
rect 36822 70694 67234 70746
rect 67286 70694 67298 70746
rect 67350 70694 67362 70746
rect 67414 70694 67426 70746
rect 67478 70694 67490 70746
rect 67542 70694 77924 70746
rect 2024 70672 77924 70694
rect 2024 70202 77924 70224
rect 2024 70150 5134 70202
rect 5186 70150 5198 70202
rect 5250 70150 5262 70202
rect 5314 70150 5326 70202
rect 5378 70150 5390 70202
rect 5442 70150 35854 70202
rect 35906 70150 35918 70202
rect 35970 70150 35982 70202
rect 36034 70150 36046 70202
rect 36098 70150 36110 70202
rect 36162 70150 66574 70202
rect 66626 70150 66638 70202
rect 66690 70150 66702 70202
rect 66754 70150 66766 70202
rect 66818 70150 66830 70202
rect 66882 70150 77924 70202
rect 2024 70128 77924 70150
rect 2024 69658 77924 69680
rect 2024 69606 5794 69658
rect 5846 69606 5858 69658
rect 5910 69606 5922 69658
rect 5974 69606 5986 69658
rect 6038 69606 6050 69658
rect 6102 69606 36514 69658
rect 36566 69606 36578 69658
rect 36630 69606 36642 69658
rect 36694 69606 36706 69658
rect 36758 69606 36770 69658
rect 36822 69606 67234 69658
rect 67286 69606 67298 69658
rect 67350 69606 67362 69658
rect 67414 69606 67426 69658
rect 67478 69606 67490 69658
rect 67542 69606 77924 69658
rect 2024 69584 77924 69606
rect 2024 69114 77924 69136
rect 2024 69062 5134 69114
rect 5186 69062 5198 69114
rect 5250 69062 5262 69114
rect 5314 69062 5326 69114
rect 5378 69062 5390 69114
rect 5442 69062 35854 69114
rect 35906 69062 35918 69114
rect 35970 69062 35982 69114
rect 36034 69062 36046 69114
rect 36098 69062 36110 69114
rect 36162 69062 66574 69114
rect 66626 69062 66638 69114
rect 66690 69062 66702 69114
rect 66754 69062 66766 69114
rect 66818 69062 66830 69114
rect 66882 69062 77924 69114
rect 2024 69040 77924 69062
rect 2024 68570 77924 68592
rect 2024 68518 5794 68570
rect 5846 68518 5858 68570
rect 5910 68518 5922 68570
rect 5974 68518 5986 68570
rect 6038 68518 6050 68570
rect 6102 68518 36514 68570
rect 36566 68518 36578 68570
rect 36630 68518 36642 68570
rect 36694 68518 36706 68570
rect 36758 68518 36770 68570
rect 36822 68518 67234 68570
rect 67286 68518 67298 68570
rect 67350 68518 67362 68570
rect 67414 68518 67426 68570
rect 67478 68518 67490 68570
rect 67542 68518 77924 68570
rect 2024 68496 77924 68518
rect 2024 68026 77924 68048
rect 2024 67974 5134 68026
rect 5186 67974 5198 68026
rect 5250 67974 5262 68026
rect 5314 67974 5326 68026
rect 5378 67974 5390 68026
rect 5442 67974 35854 68026
rect 35906 67974 35918 68026
rect 35970 67974 35982 68026
rect 36034 67974 36046 68026
rect 36098 67974 36110 68026
rect 36162 67974 66574 68026
rect 66626 67974 66638 68026
rect 66690 67974 66702 68026
rect 66754 67974 66766 68026
rect 66818 67974 66830 68026
rect 66882 67974 77924 68026
rect 2024 67952 77924 67974
rect 2024 67482 77924 67504
rect 2024 67430 5794 67482
rect 5846 67430 5858 67482
rect 5910 67430 5922 67482
rect 5974 67430 5986 67482
rect 6038 67430 6050 67482
rect 6102 67430 36514 67482
rect 36566 67430 36578 67482
rect 36630 67430 36642 67482
rect 36694 67430 36706 67482
rect 36758 67430 36770 67482
rect 36822 67430 67234 67482
rect 67286 67430 67298 67482
rect 67350 67430 67362 67482
rect 67414 67430 67426 67482
rect 67478 67430 67490 67482
rect 67542 67430 77924 67482
rect 2024 67408 77924 67430
rect 2024 66938 77924 66960
rect 2024 66886 5134 66938
rect 5186 66886 5198 66938
rect 5250 66886 5262 66938
rect 5314 66886 5326 66938
rect 5378 66886 5390 66938
rect 5442 66886 35854 66938
rect 35906 66886 35918 66938
rect 35970 66886 35982 66938
rect 36034 66886 36046 66938
rect 36098 66886 36110 66938
rect 36162 66886 66574 66938
rect 66626 66886 66638 66938
rect 66690 66886 66702 66938
rect 66754 66886 66766 66938
rect 66818 66886 66830 66938
rect 66882 66886 77924 66938
rect 2024 66864 77924 66886
rect 2024 66394 77924 66416
rect 2024 66342 5794 66394
rect 5846 66342 5858 66394
rect 5910 66342 5922 66394
rect 5974 66342 5986 66394
rect 6038 66342 6050 66394
rect 6102 66342 36514 66394
rect 36566 66342 36578 66394
rect 36630 66342 36642 66394
rect 36694 66342 36706 66394
rect 36758 66342 36770 66394
rect 36822 66342 67234 66394
rect 67286 66342 67298 66394
rect 67350 66342 67362 66394
rect 67414 66342 67426 66394
rect 67478 66342 67490 66394
rect 67542 66342 77924 66394
rect 2024 66320 77924 66342
rect 2024 65850 77924 65872
rect 2024 65798 5134 65850
rect 5186 65798 5198 65850
rect 5250 65798 5262 65850
rect 5314 65798 5326 65850
rect 5378 65798 5390 65850
rect 5442 65798 35854 65850
rect 35906 65798 35918 65850
rect 35970 65798 35982 65850
rect 36034 65798 36046 65850
rect 36098 65798 36110 65850
rect 36162 65798 66574 65850
rect 66626 65798 66638 65850
rect 66690 65798 66702 65850
rect 66754 65798 66766 65850
rect 66818 65798 66830 65850
rect 66882 65798 77924 65850
rect 2024 65776 77924 65798
rect 2024 65306 77924 65328
rect 2024 65254 5794 65306
rect 5846 65254 5858 65306
rect 5910 65254 5922 65306
rect 5974 65254 5986 65306
rect 6038 65254 6050 65306
rect 6102 65254 36514 65306
rect 36566 65254 36578 65306
rect 36630 65254 36642 65306
rect 36694 65254 36706 65306
rect 36758 65254 36770 65306
rect 36822 65254 67234 65306
rect 67286 65254 67298 65306
rect 67350 65254 67362 65306
rect 67414 65254 67426 65306
rect 67478 65254 67490 65306
rect 67542 65254 77924 65306
rect 2024 65232 77924 65254
rect 2024 64762 77924 64784
rect 2024 64710 5134 64762
rect 5186 64710 5198 64762
rect 5250 64710 5262 64762
rect 5314 64710 5326 64762
rect 5378 64710 5390 64762
rect 5442 64710 35854 64762
rect 35906 64710 35918 64762
rect 35970 64710 35982 64762
rect 36034 64710 36046 64762
rect 36098 64710 36110 64762
rect 36162 64710 66574 64762
rect 66626 64710 66638 64762
rect 66690 64710 66702 64762
rect 66754 64710 66766 64762
rect 66818 64710 66830 64762
rect 66882 64710 77924 64762
rect 2024 64688 77924 64710
rect 2024 64218 77924 64240
rect 2024 64166 5794 64218
rect 5846 64166 5858 64218
rect 5910 64166 5922 64218
rect 5974 64166 5986 64218
rect 6038 64166 6050 64218
rect 6102 64166 36514 64218
rect 36566 64166 36578 64218
rect 36630 64166 36642 64218
rect 36694 64166 36706 64218
rect 36758 64166 36770 64218
rect 36822 64166 67234 64218
rect 67286 64166 67298 64218
rect 67350 64166 67362 64218
rect 67414 64166 67426 64218
rect 67478 64166 67490 64218
rect 67542 64166 77924 64218
rect 2024 64144 77924 64166
rect 2024 63674 77924 63696
rect 2024 63622 5134 63674
rect 5186 63622 5198 63674
rect 5250 63622 5262 63674
rect 5314 63622 5326 63674
rect 5378 63622 5390 63674
rect 5442 63622 35854 63674
rect 35906 63622 35918 63674
rect 35970 63622 35982 63674
rect 36034 63622 36046 63674
rect 36098 63622 36110 63674
rect 36162 63622 66574 63674
rect 66626 63622 66638 63674
rect 66690 63622 66702 63674
rect 66754 63622 66766 63674
rect 66818 63622 66830 63674
rect 66882 63622 77924 63674
rect 2024 63600 77924 63622
rect 2024 63130 77924 63152
rect 2024 63078 5794 63130
rect 5846 63078 5858 63130
rect 5910 63078 5922 63130
rect 5974 63078 5986 63130
rect 6038 63078 6050 63130
rect 6102 63078 36514 63130
rect 36566 63078 36578 63130
rect 36630 63078 36642 63130
rect 36694 63078 36706 63130
rect 36758 63078 36770 63130
rect 36822 63078 67234 63130
rect 67286 63078 67298 63130
rect 67350 63078 67362 63130
rect 67414 63078 67426 63130
rect 67478 63078 67490 63130
rect 67542 63078 77924 63130
rect 2024 63056 77924 63078
rect 2024 62586 77924 62608
rect 2024 62534 5134 62586
rect 5186 62534 5198 62586
rect 5250 62534 5262 62586
rect 5314 62534 5326 62586
rect 5378 62534 5390 62586
rect 5442 62534 35854 62586
rect 35906 62534 35918 62586
rect 35970 62534 35982 62586
rect 36034 62534 36046 62586
rect 36098 62534 36110 62586
rect 36162 62534 66574 62586
rect 66626 62534 66638 62586
rect 66690 62534 66702 62586
rect 66754 62534 66766 62586
rect 66818 62534 66830 62586
rect 66882 62534 77924 62586
rect 2024 62512 77924 62534
rect 2024 62042 77924 62064
rect 2024 61990 5794 62042
rect 5846 61990 5858 62042
rect 5910 61990 5922 62042
rect 5974 61990 5986 62042
rect 6038 61990 6050 62042
rect 6102 61990 36514 62042
rect 36566 61990 36578 62042
rect 36630 61990 36642 62042
rect 36694 61990 36706 62042
rect 36758 61990 36770 62042
rect 36822 61990 67234 62042
rect 67286 61990 67298 62042
rect 67350 61990 67362 62042
rect 67414 61990 67426 62042
rect 67478 61990 67490 62042
rect 67542 61990 77924 62042
rect 2024 61968 77924 61990
rect 2024 61498 77924 61520
rect 2024 61446 5134 61498
rect 5186 61446 5198 61498
rect 5250 61446 5262 61498
rect 5314 61446 5326 61498
rect 5378 61446 5390 61498
rect 5442 61446 35854 61498
rect 35906 61446 35918 61498
rect 35970 61446 35982 61498
rect 36034 61446 36046 61498
rect 36098 61446 36110 61498
rect 36162 61446 66574 61498
rect 66626 61446 66638 61498
rect 66690 61446 66702 61498
rect 66754 61446 66766 61498
rect 66818 61446 66830 61498
rect 66882 61446 77924 61498
rect 2024 61424 77924 61446
rect 2024 60954 77924 60976
rect 2024 60902 5794 60954
rect 5846 60902 5858 60954
rect 5910 60902 5922 60954
rect 5974 60902 5986 60954
rect 6038 60902 6050 60954
rect 6102 60902 36514 60954
rect 36566 60902 36578 60954
rect 36630 60902 36642 60954
rect 36694 60902 36706 60954
rect 36758 60902 36770 60954
rect 36822 60902 67234 60954
rect 67286 60902 67298 60954
rect 67350 60902 67362 60954
rect 67414 60902 67426 60954
rect 67478 60902 67490 60954
rect 67542 60902 77924 60954
rect 2024 60880 77924 60902
rect 2024 60410 77924 60432
rect 2024 60358 5134 60410
rect 5186 60358 5198 60410
rect 5250 60358 5262 60410
rect 5314 60358 5326 60410
rect 5378 60358 5390 60410
rect 5442 60358 35854 60410
rect 35906 60358 35918 60410
rect 35970 60358 35982 60410
rect 36034 60358 36046 60410
rect 36098 60358 36110 60410
rect 36162 60358 66574 60410
rect 66626 60358 66638 60410
rect 66690 60358 66702 60410
rect 66754 60358 66766 60410
rect 66818 60358 66830 60410
rect 66882 60358 77924 60410
rect 2024 60336 77924 60358
rect 2024 59866 77924 59888
rect 2024 59814 5794 59866
rect 5846 59814 5858 59866
rect 5910 59814 5922 59866
rect 5974 59814 5986 59866
rect 6038 59814 6050 59866
rect 6102 59814 36514 59866
rect 36566 59814 36578 59866
rect 36630 59814 36642 59866
rect 36694 59814 36706 59866
rect 36758 59814 36770 59866
rect 36822 59814 67234 59866
rect 67286 59814 67298 59866
rect 67350 59814 67362 59866
rect 67414 59814 67426 59866
rect 67478 59814 67490 59866
rect 67542 59814 77924 59866
rect 2024 59792 77924 59814
rect 2024 59322 77924 59344
rect 2024 59270 5134 59322
rect 5186 59270 5198 59322
rect 5250 59270 5262 59322
rect 5314 59270 5326 59322
rect 5378 59270 5390 59322
rect 5442 59270 35854 59322
rect 35906 59270 35918 59322
rect 35970 59270 35982 59322
rect 36034 59270 36046 59322
rect 36098 59270 36110 59322
rect 36162 59270 66574 59322
rect 66626 59270 66638 59322
rect 66690 59270 66702 59322
rect 66754 59270 66766 59322
rect 66818 59270 66830 59322
rect 66882 59270 77924 59322
rect 2024 59248 77924 59270
rect 2024 58778 77924 58800
rect 2024 58726 5794 58778
rect 5846 58726 5858 58778
rect 5910 58726 5922 58778
rect 5974 58726 5986 58778
rect 6038 58726 6050 58778
rect 6102 58726 36514 58778
rect 36566 58726 36578 58778
rect 36630 58726 36642 58778
rect 36694 58726 36706 58778
rect 36758 58726 36770 58778
rect 36822 58726 67234 58778
rect 67286 58726 67298 58778
rect 67350 58726 67362 58778
rect 67414 58726 67426 58778
rect 67478 58726 67490 58778
rect 67542 58726 77924 58778
rect 2024 58704 77924 58726
rect 2024 58234 77924 58256
rect 2024 58182 5134 58234
rect 5186 58182 5198 58234
rect 5250 58182 5262 58234
rect 5314 58182 5326 58234
rect 5378 58182 5390 58234
rect 5442 58182 35854 58234
rect 35906 58182 35918 58234
rect 35970 58182 35982 58234
rect 36034 58182 36046 58234
rect 36098 58182 36110 58234
rect 36162 58182 66574 58234
rect 66626 58182 66638 58234
rect 66690 58182 66702 58234
rect 66754 58182 66766 58234
rect 66818 58182 66830 58234
rect 66882 58182 77924 58234
rect 2024 58160 77924 58182
rect 2024 57690 77924 57712
rect 2024 57638 5794 57690
rect 5846 57638 5858 57690
rect 5910 57638 5922 57690
rect 5974 57638 5986 57690
rect 6038 57638 6050 57690
rect 6102 57638 36514 57690
rect 36566 57638 36578 57690
rect 36630 57638 36642 57690
rect 36694 57638 36706 57690
rect 36758 57638 36770 57690
rect 36822 57638 67234 57690
rect 67286 57638 67298 57690
rect 67350 57638 67362 57690
rect 67414 57638 67426 57690
rect 67478 57638 67490 57690
rect 67542 57638 77924 57690
rect 2024 57616 77924 57638
rect 2024 57146 77924 57168
rect 2024 57094 5134 57146
rect 5186 57094 5198 57146
rect 5250 57094 5262 57146
rect 5314 57094 5326 57146
rect 5378 57094 5390 57146
rect 5442 57094 35854 57146
rect 35906 57094 35918 57146
rect 35970 57094 35982 57146
rect 36034 57094 36046 57146
rect 36098 57094 36110 57146
rect 36162 57094 66574 57146
rect 66626 57094 66638 57146
rect 66690 57094 66702 57146
rect 66754 57094 66766 57146
rect 66818 57094 66830 57146
rect 66882 57094 77924 57146
rect 2024 57072 77924 57094
rect 2024 56602 77924 56624
rect 2024 56550 5794 56602
rect 5846 56550 5858 56602
rect 5910 56550 5922 56602
rect 5974 56550 5986 56602
rect 6038 56550 6050 56602
rect 6102 56550 36514 56602
rect 36566 56550 36578 56602
rect 36630 56550 36642 56602
rect 36694 56550 36706 56602
rect 36758 56550 36770 56602
rect 36822 56550 67234 56602
rect 67286 56550 67298 56602
rect 67350 56550 67362 56602
rect 67414 56550 67426 56602
rect 67478 56550 67490 56602
rect 67542 56550 77924 56602
rect 2024 56528 77924 56550
rect 2024 56058 77924 56080
rect 2024 56006 5134 56058
rect 5186 56006 5198 56058
rect 5250 56006 5262 56058
rect 5314 56006 5326 56058
rect 5378 56006 5390 56058
rect 5442 56006 35854 56058
rect 35906 56006 35918 56058
rect 35970 56006 35982 56058
rect 36034 56006 36046 56058
rect 36098 56006 36110 56058
rect 36162 56006 66574 56058
rect 66626 56006 66638 56058
rect 66690 56006 66702 56058
rect 66754 56006 66766 56058
rect 66818 56006 66830 56058
rect 66882 56006 77924 56058
rect 2024 55984 77924 56006
rect 2024 55514 77924 55536
rect 2024 55462 5794 55514
rect 5846 55462 5858 55514
rect 5910 55462 5922 55514
rect 5974 55462 5986 55514
rect 6038 55462 6050 55514
rect 6102 55462 36514 55514
rect 36566 55462 36578 55514
rect 36630 55462 36642 55514
rect 36694 55462 36706 55514
rect 36758 55462 36770 55514
rect 36822 55462 67234 55514
rect 67286 55462 67298 55514
rect 67350 55462 67362 55514
rect 67414 55462 67426 55514
rect 67478 55462 67490 55514
rect 67542 55462 77924 55514
rect 2024 55440 77924 55462
rect 2024 54970 77924 54992
rect 2024 54918 5134 54970
rect 5186 54918 5198 54970
rect 5250 54918 5262 54970
rect 5314 54918 5326 54970
rect 5378 54918 5390 54970
rect 5442 54918 35854 54970
rect 35906 54918 35918 54970
rect 35970 54918 35982 54970
rect 36034 54918 36046 54970
rect 36098 54918 36110 54970
rect 36162 54918 66574 54970
rect 66626 54918 66638 54970
rect 66690 54918 66702 54970
rect 66754 54918 66766 54970
rect 66818 54918 66830 54970
rect 66882 54918 77924 54970
rect 2024 54896 77924 54918
rect 2024 54426 77924 54448
rect 2024 54374 5794 54426
rect 5846 54374 5858 54426
rect 5910 54374 5922 54426
rect 5974 54374 5986 54426
rect 6038 54374 6050 54426
rect 6102 54374 36514 54426
rect 36566 54374 36578 54426
rect 36630 54374 36642 54426
rect 36694 54374 36706 54426
rect 36758 54374 36770 54426
rect 36822 54374 67234 54426
rect 67286 54374 67298 54426
rect 67350 54374 67362 54426
rect 67414 54374 67426 54426
rect 67478 54374 67490 54426
rect 67542 54374 77924 54426
rect 2024 54352 77924 54374
rect 2024 53882 77924 53904
rect 2024 53830 5134 53882
rect 5186 53830 5198 53882
rect 5250 53830 5262 53882
rect 5314 53830 5326 53882
rect 5378 53830 5390 53882
rect 5442 53830 35854 53882
rect 35906 53830 35918 53882
rect 35970 53830 35982 53882
rect 36034 53830 36046 53882
rect 36098 53830 36110 53882
rect 36162 53830 66574 53882
rect 66626 53830 66638 53882
rect 66690 53830 66702 53882
rect 66754 53830 66766 53882
rect 66818 53830 66830 53882
rect 66882 53830 77924 53882
rect 2024 53808 77924 53830
rect 2024 53338 77924 53360
rect 2024 53286 5794 53338
rect 5846 53286 5858 53338
rect 5910 53286 5922 53338
rect 5974 53286 5986 53338
rect 6038 53286 6050 53338
rect 6102 53286 36514 53338
rect 36566 53286 36578 53338
rect 36630 53286 36642 53338
rect 36694 53286 36706 53338
rect 36758 53286 36770 53338
rect 36822 53286 67234 53338
rect 67286 53286 67298 53338
rect 67350 53286 67362 53338
rect 67414 53286 67426 53338
rect 67478 53286 67490 53338
rect 67542 53286 77924 53338
rect 2024 53264 77924 53286
rect 2024 52794 77924 52816
rect 2024 52742 5134 52794
rect 5186 52742 5198 52794
rect 5250 52742 5262 52794
rect 5314 52742 5326 52794
rect 5378 52742 5390 52794
rect 5442 52742 35854 52794
rect 35906 52742 35918 52794
rect 35970 52742 35982 52794
rect 36034 52742 36046 52794
rect 36098 52742 36110 52794
rect 36162 52742 66574 52794
rect 66626 52742 66638 52794
rect 66690 52742 66702 52794
rect 66754 52742 66766 52794
rect 66818 52742 66830 52794
rect 66882 52742 77924 52794
rect 2024 52720 77924 52742
rect 2024 52250 77924 52272
rect 2024 52198 5794 52250
rect 5846 52198 5858 52250
rect 5910 52198 5922 52250
rect 5974 52198 5986 52250
rect 6038 52198 6050 52250
rect 6102 52198 36514 52250
rect 36566 52198 36578 52250
rect 36630 52198 36642 52250
rect 36694 52198 36706 52250
rect 36758 52198 36770 52250
rect 36822 52198 67234 52250
rect 67286 52198 67298 52250
rect 67350 52198 67362 52250
rect 67414 52198 67426 52250
rect 67478 52198 67490 52250
rect 67542 52198 77924 52250
rect 2024 52176 77924 52198
rect 77570 51756 77576 51808
rect 77628 51756 77634 51808
rect 2024 51706 77924 51728
rect 2024 51654 5134 51706
rect 5186 51654 5198 51706
rect 5250 51654 5262 51706
rect 5314 51654 5326 51706
rect 5378 51654 5390 51706
rect 5442 51654 35854 51706
rect 35906 51654 35918 51706
rect 35970 51654 35982 51706
rect 36034 51654 36046 51706
rect 36098 51654 36110 51706
rect 36162 51654 66574 51706
rect 66626 51654 66638 51706
rect 66690 51654 66702 51706
rect 66754 51654 66766 51706
rect 66818 51654 66830 51706
rect 66882 51654 77924 51706
rect 2024 51632 77924 51654
rect 2024 51162 77924 51184
rect 2024 51110 5794 51162
rect 5846 51110 5858 51162
rect 5910 51110 5922 51162
rect 5974 51110 5986 51162
rect 6038 51110 6050 51162
rect 6102 51110 36514 51162
rect 36566 51110 36578 51162
rect 36630 51110 36642 51162
rect 36694 51110 36706 51162
rect 36758 51110 36770 51162
rect 36822 51110 67234 51162
rect 67286 51110 67298 51162
rect 67350 51110 67362 51162
rect 67414 51110 67426 51162
rect 67478 51110 67490 51162
rect 67542 51110 77924 51162
rect 2024 51088 77924 51110
rect 2024 50618 77924 50640
rect 2024 50566 5134 50618
rect 5186 50566 5198 50618
rect 5250 50566 5262 50618
rect 5314 50566 5326 50618
rect 5378 50566 5390 50618
rect 5442 50566 35854 50618
rect 35906 50566 35918 50618
rect 35970 50566 35982 50618
rect 36034 50566 36046 50618
rect 36098 50566 36110 50618
rect 36162 50566 66574 50618
rect 66626 50566 66638 50618
rect 66690 50566 66702 50618
rect 66754 50566 66766 50618
rect 66818 50566 66830 50618
rect 66882 50566 77924 50618
rect 2024 50544 77924 50566
rect 2024 50074 77924 50096
rect 2024 50022 5794 50074
rect 5846 50022 5858 50074
rect 5910 50022 5922 50074
rect 5974 50022 5986 50074
rect 6038 50022 6050 50074
rect 6102 50022 36514 50074
rect 36566 50022 36578 50074
rect 36630 50022 36642 50074
rect 36694 50022 36706 50074
rect 36758 50022 36770 50074
rect 36822 50022 67234 50074
rect 67286 50022 67298 50074
rect 67350 50022 67362 50074
rect 67414 50022 67426 50074
rect 67478 50022 67490 50074
rect 67542 50022 77924 50074
rect 2024 50000 77924 50022
rect 77570 49716 77576 49768
rect 77628 49716 77634 49768
rect 2024 49530 77924 49552
rect 2024 49478 5134 49530
rect 5186 49478 5198 49530
rect 5250 49478 5262 49530
rect 5314 49478 5326 49530
rect 5378 49478 5390 49530
rect 5442 49478 35854 49530
rect 35906 49478 35918 49530
rect 35970 49478 35982 49530
rect 36034 49478 36046 49530
rect 36098 49478 36110 49530
rect 36162 49478 66574 49530
rect 66626 49478 66638 49530
rect 66690 49478 66702 49530
rect 66754 49478 66766 49530
rect 66818 49478 66830 49530
rect 66882 49478 77924 49530
rect 2024 49456 77924 49478
rect 2024 48986 77924 49008
rect 2024 48934 5794 48986
rect 5846 48934 5858 48986
rect 5910 48934 5922 48986
rect 5974 48934 5986 48986
rect 6038 48934 6050 48986
rect 6102 48934 36514 48986
rect 36566 48934 36578 48986
rect 36630 48934 36642 48986
rect 36694 48934 36706 48986
rect 36758 48934 36770 48986
rect 36822 48934 67234 48986
rect 67286 48934 67298 48986
rect 67350 48934 67362 48986
rect 67414 48934 67426 48986
rect 67478 48934 67490 48986
rect 67542 48934 77924 48986
rect 2024 48912 77924 48934
rect 2024 48442 77924 48464
rect 2024 48390 5134 48442
rect 5186 48390 5198 48442
rect 5250 48390 5262 48442
rect 5314 48390 5326 48442
rect 5378 48390 5390 48442
rect 5442 48390 35854 48442
rect 35906 48390 35918 48442
rect 35970 48390 35982 48442
rect 36034 48390 36046 48442
rect 36098 48390 36110 48442
rect 36162 48390 66574 48442
rect 66626 48390 66638 48442
rect 66690 48390 66702 48442
rect 66754 48390 66766 48442
rect 66818 48390 66830 48442
rect 66882 48390 77924 48442
rect 2024 48368 77924 48390
rect 2024 47898 77924 47920
rect 2024 47846 5794 47898
rect 5846 47846 5858 47898
rect 5910 47846 5922 47898
rect 5974 47846 5986 47898
rect 6038 47846 6050 47898
rect 6102 47846 36514 47898
rect 36566 47846 36578 47898
rect 36630 47846 36642 47898
rect 36694 47846 36706 47898
rect 36758 47846 36770 47898
rect 36822 47846 67234 47898
rect 67286 47846 67298 47898
rect 67350 47846 67362 47898
rect 67414 47846 67426 47898
rect 67478 47846 67490 47898
rect 67542 47846 77924 47898
rect 2024 47824 77924 47846
rect 2024 47354 77924 47376
rect 2024 47302 5134 47354
rect 5186 47302 5198 47354
rect 5250 47302 5262 47354
rect 5314 47302 5326 47354
rect 5378 47302 5390 47354
rect 5442 47302 35854 47354
rect 35906 47302 35918 47354
rect 35970 47302 35982 47354
rect 36034 47302 36046 47354
rect 36098 47302 36110 47354
rect 36162 47302 66574 47354
rect 66626 47302 66638 47354
rect 66690 47302 66702 47354
rect 66754 47302 66766 47354
rect 66818 47302 66830 47354
rect 66882 47302 77924 47354
rect 2024 47280 77924 47302
rect 2024 46810 77924 46832
rect 2024 46758 5794 46810
rect 5846 46758 5858 46810
rect 5910 46758 5922 46810
rect 5974 46758 5986 46810
rect 6038 46758 6050 46810
rect 6102 46758 36514 46810
rect 36566 46758 36578 46810
rect 36630 46758 36642 46810
rect 36694 46758 36706 46810
rect 36758 46758 36770 46810
rect 36822 46758 67234 46810
rect 67286 46758 67298 46810
rect 67350 46758 67362 46810
rect 67414 46758 67426 46810
rect 67478 46758 67490 46810
rect 67542 46758 77924 46810
rect 2024 46736 77924 46758
rect 2024 46266 77924 46288
rect 2024 46214 5134 46266
rect 5186 46214 5198 46266
rect 5250 46214 5262 46266
rect 5314 46214 5326 46266
rect 5378 46214 5390 46266
rect 5442 46214 35854 46266
rect 35906 46214 35918 46266
rect 35970 46214 35982 46266
rect 36034 46214 36046 46266
rect 36098 46214 36110 46266
rect 36162 46214 66574 46266
rect 66626 46214 66638 46266
rect 66690 46214 66702 46266
rect 66754 46214 66766 46266
rect 66818 46214 66830 46266
rect 66882 46214 77924 46266
rect 2024 46192 77924 46214
rect 2024 45722 77924 45744
rect 2024 45670 5794 45722
rect 5846 45670 5858 45722
rect 5910 45670 5922 45722
rect 5974 45670 5986 45722
rect 6038 45670 6050 45722
rect 6102 45670 36514 45722
rect 36566 45670 36578 45722
rect 36630 45670 36642 45722
rect 36694 45670 36706 45722
rect 36758 45670 36770 45722
rect 36822 45670 67234 45722
rect 67286 45670 67298 45722
rect 67350 45670 67362 45722
rect 67414 45670 67426 45722
rect 67478 45670 67490 45722
rect 67542 45670 77924 45722
rect 2024 45648 77924 45670
rect 2024 45178 77924 45200
rect 2024 45126 5134 45178
rect 5186 45126 5198 45178
rect 5250 45126 5262 45178
rect 5314 45126 5326 45178
rect 5378 45126 5390 45178
rect 5442 45126 35854 45178
rect 35906 45126 35918 45178
rect 35970 45126 35982 45178
rect 36034 45126 36046 45178
rect 36098 45126 36110 45178
rect 36162 45126 66574 45178
rect 66626 45126 66638 45178
rect 66690 45126 66702 45178
rect 66754 45126 66766 45178
rect 66818 45126 66830 45178
rect 66882 45126 77924 45178
rect 2024 45104 77924 45126
rect 2024 44634 77924 44656
rect 2024 44582 5794 44634
rect 5846 44582 5858 44634
rect 5910 44582 5922 44634
rect 5974 44582 5986 44634
rect 6038 44582 6050 44634
rect 6102 44582 36514 44634
rect 36566 44582 36578 44634
rect 36630 44582 36642 44634
rect 36694 44582 36706 44634
rect 36758 44582 36770 44634
rect 36822 44582 67234 44634
rect 67286 44582 67298 44634
rect 67350 44582 67362 44634
rect 67414 44582 67426 44634
rect 67478 44582 67490 44634
rect 67542 44582 77924 44634
rect 2024 44560 77924 44582
rect 2024 44090 77924 44112
rect 2024 44038 5134 44090
rect 5186 44038 5198 44090
rect 5250 44038 5262 44090
rect 5314 44038 5326 44090
rect 5378 44038 5390 44090
rect 5442 44038 35854 44090
rect 35906 44038 35918 44090
rect 35970 44038 35982 44090
rect 36034 44038 36046 44090
rect 36098 44038 36110 44090
rect 36162 44038 66574 44090
rect 66626 44038 66638 44090
rect 66690 44038 66702 44090
rect 66754 44038 66766 44090
rect 66818 44038 66830 44090
rect 66882 44038 77924 44090
rect 2024 44016 77924 44038
rect 64874 43800 64880 43852
rect 64932 43800 64938 43852
rect 64969 43775 65027 43781
rect 64969 43741 64981 43775
rect 65015 43772 65027 43775
rect 66533 43775 66591 43781
rect 66533 43772 66545 43775
rect 65015 43744 66545 43772
rect 65015 43741 65027 43744
rect 64969 43735 65027 43741
rect 66533 43741 66545 43744
rect 66579 43741 66591 43775
rect 66533 43735 66591 43741
rect 66898 43732 66904 43784
rect 66956 43772 66962 43784
rect 67085 43775 67143 43781
rect 67085 43772 67097 43775
rect 66956 43744 67097 43772
rect 66956 43732 66962 43744
rect 67085 43741 67097 43744
rect 67131 43741 67143 43775
rect 67085 43735 67143 43741
rect 65337 43639 65395 43645
rect 65337 43605 65349 43639
rect 65383 43636 65395 43639
rect 65426 43636 65432 43648
rect 65383 43608 65432 43636
rect 65383 43605 65395 43608
rect 65337 43599 65395 43605
rect 65426 43596 65432 43608
rect 65484 43596 65490 43648
rect 2024 43546 77924 43568
rect 2024 43494 5794 43546
rect 5846 43494 5858 43546
rect 5910 43494 5922 43546
rect 5974 43494 5986 43546
rect 6038 43494 6050 43546
rect 6102 43494 36514 43546
rect 36566 43494 36578 43546
rect 36630 43494 36642 43546
rect 36694 43494 36706 43546
rect 36758 43494 36770 43546
rect 36822 43494 67234 43546
rect 67286 43494 67298 43546
rect 67350 43494 67362 43546
rect 67414 43494 67426 43546
rect 67478 43494 67490 43546
rect 67542 43494 77924 43546
rect 2024 43472 77924 43494
rect 66254 43392 66260 43444
rect 66312 43432 66318 43444
rect 66898 43432 66904 43444
rect 66312 43404 66904 43432
rect 66312 43392 66318 43404
rect 66898 43392 66904 43404
rect 66956 43392 66962 43444
rect 65426 43324 65432 43376
rect 65484 43324 65490 43376
rect 67085 43367 67143 43373
rect 67085 43364 67097 43367
rect 66654 43336 67097 43364
rect 67085 43333 67097 43336
rect 67131 43333 67143 43367
rect 67085 43327 67143 43333
rect 67177 43299 67235 43305
rect 67177 43296 67189 43299
rect 67100 43268 67189 43296
rect 67100 43240 67128 43268
rect 67177 43265 67189 43268
rect 67223 43265 67235 43299
rect 67177 43259 67235 43265
rect 65150 43188 65156 43240
rect 65208 43188 65214 43240
rect 67082 43188 67088 43240
rect 67140 43188 67146 43240
rect 2024 43002 77924 43024
rect 2024 42950 5134 43002
rect 5186 42950 5198 43002
rect 5250 42950 5262 43002
rect 5314 42950 5326 43002
rect 5378 42950 5390 43002
rect 5442 42950 35854 43002
rect 35906 42950 35918 43002
rect 35970 42950 35982 43002
rect 36034 42950 36046 43002
rect 36098 42950 36110 43002
rect 36162 42950 66574 43002
rect 66626 42950 66638 43002
rect 66690 42950 66702 43002
rect 66754 42950 66766 43002
rect 66818 42950 66830 43002
rect 66882 42950 77924 43002
rect 2024 42928 77924 42950
rect 59357 42755 59415 42761
rect 59357 42721 59369 42755
rect 59403 42752 59415 42755
rect 59998 42752 60004 42764
rect 59403 42724 60004 42752
rect 59403 42721 59415 42724
rect 59357 42715 59415 42721
rect 59998 42712 60004 42724
rect 60056 42752 60062 42764
rect 60093 42755 60151 42761
rect 60093 42752 60105 42755
rect 60056 42724 60105 42752
rect 60056 42712 60062 42724
rect 60093 42721 60105 42724
rect 60139 42721 60151 42755
rect 60093 42715 60151 42721
rect 57606 42644 57612 42696
rect 57664 42644 57670 42696
rect 57885 42619 57943 42625
rect 57885 42585 57897 42619
rect 57931 42616 57943 42619
rect 57974 42616 57980 42628
rect 57931 42588 57980 42616
rect 57931 42585 57943 42588
rect 57885 42579 57943 42585
rect 57974 42576 57980 42588
rect 58032 42576 58038 42628
rect 58894 42576 58900 42628
rect 58952 42576 58958 42628
rect 59538 42508 59544 42560
rect 59596 42508 59602 42560
rect 2024 42458 77924 42480
rect 2024 42406 5794 42458
rect 5846 42406 5858 42458
rect 5910 42406 5922 42458
rect 5974 42406 5986 42458
rect 6038 42406 6050 42458
rect 6102 42406 36514 42458
rect 36566 42406 36578 42458
rect 36630 42406 36642 42458
rect 36694 42406 36706 42458
rect 36758 42406 36770 42458
rect 36822 42406 67234 42458
rect 67286 42406 67298 42458
rect 67350 42406 67362 42458
rect 67414 42406 67426 42458
rect 67478 42406 67490 42458
rect 67542 42406 77924 42458
rect 2024 42384 77924 42406
rect 57974 42304 57980 42356
rect 58032 42344 58038 42356
rect 58069 42347 58127 42353
rect 58069 42344 58081 42347
rect 58032 42316 58081 42344
rect 58032 42304 58038 42316
rect 58069 42313 58081 42316
rect 58115 42313 58127 42347
rect 58069 42307 58127 42313
rect 58894 42304 58900 42356
rect 58952 42304 58958 42356
rect 59538 42276 59544 42288
rect 58176 42248 59544 42276
rect 58176 42217 58204 42248
rect 59538 42236 59544 42248
rect 59596 42236 59602 42288
rect 58161 42211 58219 42217
rect 58161 42177 58173 42211
rect 58207 42177 58219 42211
rect 58161 42171 58219 42177
rect 58986 42168 58992 42220
rect 59044 42168 59050 42220
rect 2024 41914 77924 41936
rect 2024 41862 5134 41914
rect 5186 41862 5198 41914
rect 5250 41862 5262 41914
rect 5314 41862 5326 41914
rect 5378 41862 5390 41914
rect 5442 41862 35854 41914
rect 35906 41862 35918 41914
rect 35970 41862 35982 41914
rect 36034 41862 36046 41914
rect 36098 41862 36110 41914
rect 36162 41862 66574 41914
rect 66626 41862 66638 41914
rect 66690 41862 66702 41914
rect 66754 41862 66766 41914
rect 66818 41862 66830 41914
rect 66882 41862 77924 41914
rect 2024 41840 77924 41862
rect 64693 41803 64751 41809
rect 64693 41769 64705 41803
rect 64739 41800 64751 41803
rect 64874 41800 64880 41812
rect 64739 41772 64880 41800
rect 64739 41769 64751 41772
rect 64693 41763 64751 41769
rect 64874 41760 64880 41772
rect 64932 41760 64938 41812
rect 71332 41636 76420 41664
rect 1210 41556 1216 41608
rect 1268 41596 1274 41608
rect 2317 41599 2375 41605
rect 2317 41596 2329 41599
rect 1268 41568 2329 41596
rect 1268 41556 1274 41568
rect 2317 41565 2329 41568
rect 2363 41565 2375 41599
rect 2317 41559 2375 41565
rect 64598 41556 64604 41608
rect 64656 41556 64662 41608
rect 64782 41556 64788 41608
rect 64840 41556 64846 41608
rect 71332 41605 71360 41636
rect 76392 41608 76420 41636
rect 71317 41599 71375 41605
rect 71317 41565 71329 41599
rect 71363 41565 71375 41599
rect 71317 41559 71375 41565
rect 74350 41556 74356 41608
rect 74408 41556 74414 41608
rect 76374 41556 76380 41608
rect 76432 41556 76438 41608
rect 74626 41488 74632 41540
rect 74684 41488 74690 41540
rect 76285 41531 76343 41537
rect 76285 41528 76297 41531
rect 75854 41500 76297 41528
rect 76285 41497 76297 41500
rect 76331 41497 76343 41531
rect 76285 41491 76343 41497
rect 71222 41420 71228 41472
rect 71280 41420 71286 41472
rect 75914 41420 75920 41472
rect 75972 41460 75978 41472
rect 76101 41463 76159 41469
rect 76101 41460 76113 41463
rect 75972 41432 76113 41460
rect 75972 41420 75978 41432
rect 76101 41429 76113 41432
rect 76147 41429 76159 41463
rect 76101 41423 76159 41429
rect 2024 41370 77924 41392
rect 2024 41318 5794 41370
rect 5846 41318 5858 41370
rect 5910 41318 5922 41370
rect 5974 41318 5986 41370
rect 6038 41318 6050 41370
rect 6102 41318 36514 41370
rect 36566 41318 36578 41370
rect 36630 41318 36642 41370
rect 36694 41318 36706 41370
rect 36758 41318 36770 41370
rect 36822 41318 67234 41370
rect 67286 41318 67298 41370
rect 67350 41318 67362 41370
rect 67414 41318 67426 41370
rect 67478 41318 67490 41370
rect 67542 41318 77924 41370
rect 2024 41296 77924 41318
rect 74350 41256 74356 41268
rect 70228 41228 74356 41256
rect 68278 41080 68284 41132
rect 68336 41120 68342 41132
rect 70228 41129 70256 41228
rect 74350 41216 74356 41228
rect 74408 41216 74414 41268
rect 71222 41148 71228 41200
rect 71280 41148 71286 41200
rect 70213 41123 70271 41129
rect 70213 41120 70225 41123
rect 68336 41092 70225 41120
rect 68336 41080 68342 41092
rect 70213 41089 70225 41092
rect 70259 41089 70271 41123
rect 70213 41083 70271 41089
rect 74445 41123 74503 41129
rect 74445 41089 74457 41123
rect 74491 41120 74503 41123
rect 75273 41123 75331 41129
rect 75273 41120 75285 41123
rect 74491 41092 75285 41120
rect 74491 41089 74503 41092
rect 74445 41083 74503 41089
rect 75273 41089 75285 41092
rect 75319 41089 75331 41123
rect 75273 41083 75331 41089
rect 70486 41012 70492 41064
rect 70544 41012 70550 41064
rect 71130 41012 71136 41064
rect 71188 41052 71194 41064
rect 74353 41055 74411 41061
rect 74353 41052 74365 41055
rect 71188 41024 74365 41052
rect 71188 41012 71194 41024
rect 74353 41021 74365 41024
rect 74399 41021 74411 41055
rect 74353 41015 74411 41021
rect 74626 41012 74632 41064
rect 74684 41052 74690 41064
rect 74813 41055 74871 41061
rect 74813 41052 74825 41055
rect 74684 41024 74825 41052
rect 74684 41012 74690 41024
rect 74813 41021 74825 41024
rect 74859 41021 74871 41055
rect 74813 41015 74871 41021
rect 75914 41012 75920 41064
rect 75972 41012 75978 41064
rect 71958 40876 71964 40928
rect 72016 40876 72022 40928
rect 2024 40826 77924 40848
rect 2024 40774 5134 40826
rect 5186 40774 5198 40826
rect 5250 40774 5262 40826
rect 5314 40774 5326 40826
rect 5378 40774 5390 40826
rect 5442 40774 35854 40826
rect 35906 40774 35918 40826
rect 35970 40774 35982 40826
rect 36034 40774 36046 40826
rect 36098 40774 36110 40826
rect 36162 40774 66574 40826
rect 66626 40774 66638 40826
rect 66690 40774 66702 40826
rect 66754 40774 66766 40826
rect 66818 40774 66830 40826
rect 66882 40774 77924 40826
rect 2024 40752 77924 40774
rect 61197 40715 61255 40721
rect 61197 40681 61209 40715
rect 61243 40712 61255 40715
rect 61638 40715 61696 40721
rect 61638 40712 61650 40715
rect 61243 40684 61650 40712
rect 61243 40681 61255 40684
rect 61197 40675 61255 40681
rect 61638 40681 61650 40684
rect 61684 40681 61696 40715
rect 61638 40675 61696 40681
rect 70486 40672 70492 40724
rect 70544 40712 70550 40724
rect 70673 40715 70731 40721
rect 70673 40712 70685 40715
rect 70544 40684 70685 40712
rect 70544 40672 70550 40684
rect 70673 40681 70685 40684
rect 70719 40681 70731 40715
rect 70673 40675 70731 40681
rect 62666 40604 62672 40656
rect 62724 40644 62730 40656
rect 63129 40647 63187 40653
rect 63129 40644 63141 40647
rect 62724 40616 63141 40644
rect 62724 40604 62730 40616
rect 63129 40613 63141 40616
rect 63175 40644 63187 40647
rect 64782 40644 64788 40656
rect 63175 40616 64788 40644
rect 63175 40613 63187 40616
rect 63129 40607 63187 40613
rect 64782 40604 64788 40616
rect 64840 40604 64846 40656
rect 66533 40647 66591 40653
rect 66533 40613 66545 40647
rect 66579 40644 66591 40647
rect 66898 40644 66904 40656
rect 66579 40616 66904 40644
rect 66579 40613 66591 40616
rect 66533 40607 66591 40613
rect 60918 40536 60924 40588
rect 60976 40536 60982 40588
rect 63494 40576 63500 40588
rect 61396 40548 63500 40576
rect 60826 40468 60832 40520
rect 60884 40468 60890 40520
rect 61396 40517 61424 40548
rect 63494 40536 63500 40548
rect 63552 40576 63558 40588
rect 65150 40576 65156 40588
rect 63552 40548 65156 40576
rect 63552 40536 63558 40548
rect 65150 40536 65156 40548
rect 65208 40536 65214 40588
rect 65889 40579 65947 40585
rect 65889 40576 65901 40579
rect 65720 40548 65901 40576
rect 61381 40511 61439 40517
rect 61381 40477 61393 40511
rect 61427 40477 61439 40511
rect 61381 40471 61439 40477
rect 57606 40400 57612 40452
rect 57664 40440 57670 40452
rect 61396 40440 61424 40471
rect 64782 40468 64788 40520
rect 64840 40508 64846 40520
rect 65720 40508 65748 40548
rect 65889 40545 65901 40548
rect 65935 40576 65947 40579
rect 66162 40576 66168 40588
rect 65935 40548 66168 40576
rect 65935 40545 65947 40548
rect 65889 40539 65947 40545
rect 66162 40536 66168 40548
rect 66220 40536 66226 40588
rect 64840 40480 65748 40508
rect 65797 40511 65855 40517
rect 64840 40468 64846 40480
rect 65797 40477 65809 40511
rect 65843 40477 65855 40511
rect 65797 40471 65855 40477
rect 57664 40412 61424 40440
rect 57664 40400 57670 40412
rect 62114 40400 62120 40452
rect 62172 40400 62178 40452
rect 65812 40440 65840 40471
rect 65978 40468 65984 40520
rect 66036 40468 66042 40520
rect 66070 40468 66076 40520
rect 66128 40468 66134 40520
rect 66548 40440 66576 40607
rect 66898 40604 66904 40616
rect 66956 40604 66962 40656
rect 70857 40647 70915 40653
rect 70857 40613 70869 40647
rect 70903 40644 70915 40647
rect 71498 40644 71504 40656
rect 70903 40616 71504 40644
rect 70903 40613 70915 40616
rect 70857 40607 70915 40613
rect 71498 40604 71504 40616
rect 71556 40604 71562 40656
rect 68278 40536 68284 40588
rect 68336 40536 68342 40588
rect 71130 40536 71136 40588
rect 71188 40536 71194 40588
rect 65812 40412 66576 40440
rect 66990 40400 66996 40452
rect 67048 40400 67054 40452
rect 68002 40400 68008 40452
rect 68060 40400 68066 40452
rect 60918 40332 60924 40384
rect 60976 40372 60982 40384
rect 64598 40372 64604 40384
rect 60976 40344 64604 40372
rect 60976 40332 60982 40344
rect 64598 40332 64604 40344
rect 64656 40332 64662 40384
rect 66257 40375 66315 40381
rect 66257 40341 66269 40375
rect 66303 40372 66315 40375
rect 66438 40372 66444 40384
rect 66303 40344 66444 40372
rect 66303 40341 66315 40344
rect 66257 40335 66315 40341
rect 66438 40332 66444 40344
rect 66496 40332 66502 40384
rect 2024 40282 77924 40304
rect 2024 40230 5794 40282
rect 5846 40230 5858 40282
rect 5910 40230 5922 40282
rect 5974 40230 5986 40282
rect 6038 40230 6050 40282
rect 6102 40230 36514 40282
rect 36566 40230 36578 40282
rect 36630 40230 36642 40282
rect 36694 40230 36706 40282
rect 36758 40230 36770 40282
rect 36822 40230 67234 40282
rect 67286 40230 67298 40282
rect 67350 40230 67362 40282
rect 67414 40230 67426 40282
rect 67478 40230 67490 40282
rect 67542 40230 77924 40282
rect 2024 40208 77924 40230
rect 60826 40128 60832 40180
rect 60884 40168 60890 40180
rect 62025 40171 62083 40177
rect 62025 40168 62037 40171
rect 60884 40140 62037 40168
rect 60884 40128 60890 40140
rect 62025 40137 62037 40140
rect 62071 40137 62083 40171
rect 62025 40131 62083 40137
rect 64598 40128 64604 40180
rect 64656 40168 64662 40180
rect 65797 40171 65855 40177
rect 65797 40168 65809 40171
rect 64656 40140 65809 40168
rect 64656 40128 64662 40140
rect 65797 40137 65809 40140
rect 65843 40168 65855 40171
rect 66070 40168 66076 40180
rect 65843 40140 66076 40168
rect 65843 40137 65855 40140
rect 65797 40131 65855 40137
rect 66070 40128 66076 40140
rect 66128 40128 66134 40180
rect 66717 40171 66775 40177
rect 66717 40137 66729 40171
rect 66763 40168 66775 40171
rect 68002 40168 68008 40180
rect 66763 40140 68008 40168
rect 66763 40137 66775 40140
rect 66717 40131 66775 40137
rect 68002 40128 68008 40140
rect 68060 40128 68066 40180
rect 65889 40103 65947 40109
rect 65889 40069 65901 40103
rect 65935 40100 65947 40103
rect 65935 40072 66116 40100
rect 65935 40069 65947 40072
rect 65889 40063 65947 40069
rect 58986 39992 58992 40044
rect 59044 40032 59050 40044
rect 61749 40035 61807 40041
rect 61749 40032 61761 40035
rect 59044 40004 61761 40032
rect 59044 39992 59050 40004
rect 61749 40001 61761 40004
rect 61795 40001 61807 40035
rect 61749 39995 61807 40001
rect 61841 40035 61899 40041
rect 61841 40001 61853 40035
rect 61887 40032 61899 40035
rect 62114 40032 62120 40044
rect 61887 40004 62120 40032
rect 61887 40001 61899 40004
rect 61841 39995 61899 40001
rect 62114 39992 62120 40004
rect 62172 39992 62178 40044
rect 62666 39992 62672 40044
rect 62724 39992 62730 40044
rect 65978 39992 65984 40044
rect 66036 39992 66042 40044
rect 66088 40032 66116 40072
rect 66162 40060 66168 40112
rect 66220 40060 66226 40112
rect 66898 40032 66904 40044
rect 66088 40004 66904 40032
rect 66898 39992 66904 40004
rect 66956 39992 66962 40044
rect 66990 39992 66996 40044
rect 67048 40032 67054 40044
rect 67177 40035 67235 40041
rect 67177 40032 67189 40035
rect 67048 40004 67189 40032
rect 67048 39992 67054 40004
rect 67177 40001 67189 40004
rect 67223 40001 67235 40035
rect 67177 39995 67235 40001
rect 67269 40035 67327 40041
rect 67269 40001 67281 40035
rect 67315 40001 67327 40035
rect 67269 39995 67327 40001
rect 66257 39967 66315 39973
rect 66257 39933 66269 39967
rect 66303 39933 66315 39967
rect 66257 39927 66315 39933
rect 65613 39831 65671 39837
rect 65613 39797 65625 39831
rect 65659 39828 65671 39831
rect 65794 39828 65800 39840
rect 65659 39800 65800 39828
rect 65659 39797 65671 39800
rect 65613 39791 65671 39797
rect 65794 39788 65800 39800
rect 65852 39828 65858 39840
rect 66272 39828 66300 39927
rect 67082 39924 67088 39976
rect 67140 39964 67146 39976
rect 67284 39964 67312 39995
rect 67140 39936 67312 39964
rect 67140 39924 67146 39936
rect 66438 39856 66444 39908
rect 66496 39896 66502 39908
rect 66533 39899 66591 39905
rect 66533 39896 66545 39899
rect 66496 39868 66545 39896
rect 66496 39856 66502 39868
rect 66533 39865 66545 39868
rect 66579 39865 66591 39899
rect 66533 39859 66591 39865
rect 65852 39800 66300 39828
rect 65852 39788 65858 39800
rect 2024 39738 77924 39760
rect 2024 39686 5134 39738
rect 5186 39686 5198 39738
rect 5250 39686 5262 39738
rect 5314 39686 5326 39738
rect 5378 39686 5390 39738
rect 5442 39686 35854 39738
rect 35906 39686 35918 39738
rect 35970 39686 35982 39738
rect 36034 39686 36046 39738
rect 36098 39686 36110 39738
rect 36162 39686 66574 39738
rect 66626 39686 66638 39738
rect 66690 39686 66702 39738
rect 66754 39686 66766 39738
rect 66818 39686 66830 39738
rect 66882 39686 77924 39738
rect 2024 39664 77924 39686
rect 70857 39627 70915 39633
rect 70857 39593 70869 39627
rect 70903 39624 70915 39627
rect 71130 39624 71136 39636
rect 70903 39596 71136 39624
rect 70903 39593 70915 39596
rect 70857 39587 70915 39593
rect 71130 39584 71136 39596
rect 71188 39584 71194 39636
rect 66162 39516 66168 39568
rect 66220 39556 66226 39568
rect 66533 39559 66591 39565
rect 66533 39556 66545 39559
rect 66220 39528 66545 39556
rect 66220 39516 66226 39528
rect 66533 39525 66545 39528
rect 66579 39525 66591 39559
rect 66533 39519 66591 39525
rect 76190 39516 76196 39568
rect 76248 39516 76254 39568
rect 56781 39491 56839 39497
rect 56781 39457 56793 39491
rect 56827 39488 56839 39491
rect 57606 39488 57612 39500
rect 56827 39460 57612 39488
rect 56827 39457 56839 39460
rect 56781 39451 56839 39457
rect 57606 39448 57612 39460
rect 57664 39448 57670 39500
rect 58342 39380 58348 39432
rect 58400 39420 58406 39432
rect 58805 39423 58863 39429
rect 58805 39420 58817 39423
rect 58400 39392 58817 39420
rect 58400 39380 58406 39392
rect 58805 39389 58817 39392
rect 58851 39420 58863 39423
rect 58986 39420 58992 39432
rect 58851 39392 58992 39420
rect 58851 39389 58863 39392
rect 58805 39383 58863 39389
rect 58986 39380 58992 39392
rect 59044 39380 59050 39432
rect 66254 39380 66260 39432
rect 66312 39420 66318 39432
rect 66717 39423 66775 39429
rect 66717 39420 66729 39423
rect 66312 39392 66729 39420
rect 66312 39380 66318 39392
rect 66717 39389 66729 39392
rect 66763 39389 66775 39423
rect 66717 39383 66775 39389
rect 66809 39423 66867 39429
rect 66809 39389 66821 39423
rect 66855 39420 66867 39423
rect 66898 39420 66904 39432
rect 66855 39392 66904 39420
rect 66855 39389 66867 39392
rect 66809 39383 66867 39389
rect 66898 39380 66904 39392
rect 66956 39380 66962 39432
rect 75730 39380 75736 39432
rect 75788 39420 75794 39432
rect 75917 39423 75975 39429
rect 75917 39420 75929 39423
rect 75788 39392 75929 39420
rect 75788 39380 75794 39392
rect 75917 39389 75929 39392
rect 75963 39389 75975 39423
rect 75917 39383 75975 39389
rect 57054 39312 57060 39364
rect 57112 39312 57118 39364
rect 58713 39355 58771 39361
rect 58713 39352 58725 39355
rect 58282 39324 58725 39352
rect 58713 39321 58725 39324
rect 58759 39321 58771 39355
rect 58713 39315 58771 39321
rect 70670 39312 70676 39364
rect 70728 39352 70734 39364
rect 71133 39355 71191 39361
rect 71133 39352 71145 39355
rect 70728 39324 71145 39352
rect 70728 39312 70734 39324
rect 71133 39321 71145 39324
rect 71179 39321 71191 39355
rect 71133 39315 71191 39321
rect 71409 39355 71467 39361
rect 71409 39321 71421 39355
rect 71455 39352 71467 39355
rect 71590 39352 71596 39364
rect 71455 39324 71596 39352
rect 71455 39321 71467 39324
rect 71409 39315 71467 39321
rect 71590 39312 71596 39324
rect 71648 39312 71654 39364
rect 75822 39312 75828 39364
rect 75880 39352 75886 39364
rect 76193 39355 76251 39361
rect 76193 39352 76205 39355
rect 75880 39324 76205 39352
rect 75880 39312 75886 39324
rect 76193 39321 76205 39324
rect 76239 39321 76251 39355
rect 76193 39315 76251 39321
rect 57974 39244 57980 39296
rect 58032 39284 58038 39296
rect 58529 39287 58587 39293
rect 58529 39284 58541 39287
rect 58032 39256 58541 39284
rect 58032 39244 58038 39256
rect 58529 39253 58541 39256
rect 58575 39253 58587 39287
rect 58529 39247 58587 39253
rect 66898 39244 66904 39296
rect 66956 39244 66962 39296
rect 67082 39244 67088 39296
rect 67140 39244 67146 39296
rect 71038 39244 71044 39296
rect 71096 39244 71102 39296
rect 71222 39244 71228 39296
rect 71280 39244 71286 39296
rect 76006 39244 76012 39296
rect 76064 39244 76070 39296
rect 2024 39194 77924 39216
rect 2024 39142 5794 39194
rect 5846 39142 5858 39194
rect 5910 39142 5922 39194
rect 5974 39142 5986 39194
rect 6038 39142 6050 39194
rect 6102 39142 36514 39194
rect 36566 39142 36578 39194
rect 36630 39142 36642 39194
rect 36694 39142 36706 39194
rect 36758 39142 36770 39194
rect 36822 39142 67234 39194
rect 67286 39142 67298 39194
rect 67350 39142 67362 39194
rect 67414 39142 67426 39194
rect 67478 39142 67490 39194
rect 67542 39142 77924 39194
rect 2024 39120 77924 39142
rect 71130 39040 71136 39092
rect 71188 39040 71194 39092
rect 71498 39040 71504 39092
rect 71556 39040 71562 39092
rect 71590 39040 71596 39092
rect 71648 39040 71654 39092
rect 75457 39083 75515 39089
rect 75457 39049 75469 39083
rect 75503 39080 75515 39083
rect 75914 39080 75920 39092
rect 75503 39052 75920 39080
rect 75503 39049 75515 39052
rect 75457 39043 75515 39049
rect 75914 39040 75920 39052
rect 75972 39040 75978 39092
rect 71792 38984 75684 39012
rect 1302 38904 1308 38956
rect 1360 38944 1366 38956
rect 65429 38947 65487 38953
rect 65429 38944 65441 38947
rect 1360 38916 65441 38944
rect 1360 38904 1366 38916
rect 65429 38913 65441 38916
rect 65475 38913 65487 38947
rect 65429 38907 65487 38913
rect 70857 38947 70915 38953
rect 70857 38913 70869 38947
rect 70903 38944 70915 38947
rect 71038 38944 71044 38956
rect 70903 38916 71044 38944
rect 70903 38913 70915 38916
rect 70857 38907 70915 38913
rect 71038 38904 71044 38916
rect 71096 38904 71102 38956
rect 71792 38953 71820 38984
rect 71225 38947 71283 38953
rect 71225 38913 71237 38947
rect 71271 38944 71283 38947
rect 71777 38947 71835 38953
rect 71777 38944 71789 38947
rect 71271 38916 71789 38944
rect 71271 38913 71283 38916
rect 71225 38907 71283 38913
rect 71777 38913 71789 38916
rect 71823 38913 71835 38947
rect 71777 38907 71835 38913
rect 71958 38904 71964 38956
rect 72016 38944 72022 38956
rect 74626 38944 74632 38956
rect 72016 38916 74632 38944
rect 72016 38904 72022 38916
rect 74626 38904 74632 38916
rect 74684 38944 74690 38956
rect 75549 38947 75607 38953
rect 75549 38944 75561 38947
rect 74684 38916 75561 38944
rect 74684 38904 74690 38916
rect 75549 38913 75561 38916
rect 75595 38913 75607 38947
rect 75549 38907 75607 38913
rect 70670 38836 70676 38888
rect 70728 38876 70734 38888
rect 70949 38879 71007 38885
rect 70949 38876 70961 38879
rect 70728 38848 70961 38876
rect 70728 38836 70734 38848
rect 70949 38845 70961 38848
rect 70995 38845 71007 38879
rect 70949 38839 71007 38845
rect 71317 38879 71375 38885
rect 71317 38845 71329 38879
rect 71363 38876 71375 38879
rect 71976 38876 72004 38904
rect 71363 38848 72004 38876
rect 75365 38879 75423 38885
rect 71363 38845 71375 38848
rect 71317 38839 71375 38845
rect 75365 38845 75377 38879
rect 75411 38876 75423 38879
rect 75656 38876 75684 38984
rect 76282 38904 76288 38956
rect 76340 38944 76346 38956
rect 77297 38947 77355 38953
rect 77297 38944 77309 38947
rect 76340 38916 77309 38944
rect 76340 38904 76346 38916
rect 77297 38913 77309 38916
rect 77343 38913 77355 38947
rect 77297 38907 77355 38913
rect 75730 38876 75736 38888
rect 75411 38848 75736 38876
rect 75411 38845 75423 38848
rect 75365 38839 75423 38845
rect 75730 38836 75736 38848
rect 75788 38836 75794 38888
rect 77478 38768 77484 38820
rect 77536 38768 77542 38820
rect 66438 38700 66444 38752
rect 66496 38740 66502 38752
rect 66717 38743 66775 38749
rect 66717 38740 66729 38743
rect 66496 38712 66729 38740
rect 66496 38700 66502 38712
rect 66717 38709 66729 38712
rect 66763 38709 66775 38743
rect 66717 38703 66775 38709
rect 75362 38700 75368 38752
rect 75420 38740 75426 38752
rect 75822 38740 75828 38752
rect 75420 38712 75828 38740
rect 75420 38700 75426 38712
rect 75822 38700 75828 38712
rect 75880 38740 75886 38752
rect 75917 38743 75975 38749
rect 75917 38740 75929 38743
rect 75880 38712 75929 38740
rect 75880 38700 75886 38712
rect 75917 38709 75929 38712
rect 75963 38709 75975 38743
rect 75917 38703 75975 38709
rect 2024 38650 77924 38672
rect 2024 38598 5134 38650
rect 5186 38598 5198 38650
rect 5250 38598 5262 38650
rect 5314 38598 5326 38650
rect 5378 38598 5390 38650
rect 5442 38598 35854 38650
rect 35906 38598 35918 38650
rect 35970 38598 35982 38650
rect 36034 38598 36046 38650
rect 36098 38598 36110 38650
rect 36162 38598 66574 38650
rect 66626 38598 66638 38650
rect 66690 38598 66702 38650
rect 66754 38598 66766 38650
rect 66818 38598 66830 38650
rect 66882 38598 77924 38650
rect 2024 38576 77924 38598
rect 57054 38496 57060 38548
rect 57112 38496 57118 38548
rect 63405 38539 63463 38545
rect 63405 38505 63417 38539
rect 63451 38536 63463 38539
rect 63494 38536 63500 38548
rect 63451 38508 63500 38536
rect 63451 38505 63463 38508
rect 63405 38499 63463 38505
rect 63494 38496 63500 38508
rect 63552 38496 63558 38548
rect 68278 38496 68284 38548
rect 68336 38536 68342 38548
rect 68922 38536 68928 38548
rect 68336 38508 68928 38536
rect 68336 38496 68342 38508
rect 68922 38496 68928 38508
rect 68980 38536 68986 38548
rect 69109 38539 69167 38545
rect 69109 38536 69121 38539
rect 68980 38508 69121 38536
rect 68980 38496 68986 38508
rect 69109 38505 69121 38508
rect 69155 38505 69167 38539
rect 69109 38499 69167 38505
rect 74721 38539 74779 38545
rect 74721 38505 74733 38539
rect 74767 38536 74779 38539
rect 76006 38536 76012 38548
rect 74767 38508 76012 38536
rect 74767 38505 74779 38508
rect 74721 38499 74779 38505
rect 76006 38496 76012 38508
rect 76064 38496 76070 38548
rect 76282 38496 76288 38548
rect 76340 38496 76346 38548
rect 57241 38335 57299 38341
rect 57241 38301 57253 38335
rect 57287 38301 57299 38335
rect 57241 38295 57299 38301
rect 57256 38264 57284 38295
rect 57330 38292 57336 38344
rect 57388 38292 57394 38344
rect 74626 38292 74632 38344
rect 74684 38292 74690 38344
rect 76098 38292 76104 38344
rect 76156 38292 76162 38344
rect 76282 38292 76288 38344
rect 76340 38332 76346 38344
rect 77297 38335 77355 38341
rect 77297 38332 77309 38335
rect 76340 38304 77309 38332
rect 76340 38292 76346 38304
rect 77297 38301 77309 38304
rect 77343 38301 77355 38335
rect 77297 38295 77355 38301
rect 57609 38267 57667 38273
rect 57609 38264 57621 38267
rect 57256 38236 57621 38264
rect 57609 38233 57621 38236
rect 57655 38233 57667 38267
rect 57609 38227 57667 38233
rect 57790 38224 57796 38276
rect 57848 38224 57854 38276
rect 57974 38224 57980 38276
rect 58032 38224 58038 38276
rect 64693 38267 64751 38273
rect 64693 38233 64705 38267
rect 64739 38264 64751 38267
rect 66438 38264 66444 38276
rect 64739 38236 66444 38264
rect 64739 38233 64751 38236
rect 64693 38227 64751 38233
rect 66438 38224 66444 38236
rect 66496 38264 66502 38276
rect 67821 38267 67879 38273
rect 67821 38264 67833 38267
rect 66496 38236 67833 38264
rect 66496 38224 66502 38236
rect 67821 38233 67833 38236
rect 67867 38233 67879 38267
rect 67821 38227 67879 38233
rect 77478 38156 77484 38208
rect 77536 38156 77542 38208
rect 2024 38106 77924 38128
rect 2024 38054 5794 38106
rect 5846 38054 5858 38106
rect 5910 38054 5922 38106
rect 5974 38054 5986 38106
rect 6038 38054 6050 38106
rect 6102 38054 36514 38106
rect 36566 38054 36578 38106
rect 36630 38054 36642 38106
rect 36694 38054 36706 38106
rect 36758 38054 36770 38106
rect 36822 38054 67234 38106
rect 67286 38054 67298 38106
rect 67350 38054 67362 38106
rect 67414 38054 67426 38106
rect 67478 38054 67490 38106
rect 67542 38054 77924 38106
rect 2024 38032 77924 38054
rect 67913 37927 67971 37933
rect 67913 37893 67925 37927
rect 67959 37924 67971 37927
rect 68278 37924 68284 37936
rect 67959 37896 68284 37924
rect 67959 37893 67971 37896
rect 67913 37887 67971 37893
rect 68278 37884 68284 37896
rect 68336 37884 68342 37936
rect 76466 37816 76472 37868
rect 76524 37856 76530 37868
rect 77297 37859 77355 37865
rect 77297 37856 77309 37859
rect 76524 37828 77309 37856
rect 76524 37816 76530 37828
rect 77297 37825 77309 37828
rect 77343 37825 77355 37859
rect 77297 37819 77355 37825
rect 77478 37612 77484 37664
rect 77536 37612 77542 37664
rect 2024 37562 77924 37584
rect 2024 37510 5134 37562
rect 5186 37510 5198 37562
rect 5250 37510 5262 37562
rect 5314 37510 5326 37562
rect 5378 37510 5390 37562
rect 5442 37510 35854 37562
rect 35906 37510 35918 37562
rect 35970 37510 35982 37562
rect 36034 37510 36046 37562
rect 36098 37510 36110 37562
rect 36162 37510 66574 37562
rect 66626 37510 66638 37562
rect 66690 37510 66702 37562
rect 66754 37510 66766 37562
rect 66818 37510 66830 37562
rect 66882 37510 77924 37562
rect 2024 37488 77924 37510
rect 63494 37272 63500 37324
rect 63552 37312 63558 37324
rect 64325 37315 64383 37321
rect 64325 37312 64337 37315
rect 63552 37284 64337 37312
rect 63552 37272 63558 37284
rect 64325 37281 64337 37284
rect 64371 37281 64383 37315
rect 64325 37275 64383 37281
rect 64601 37315 64659 37321
rect 64601 37281 64613 37315
rect 64647 37312 64659 37315
rect 65334 37312 65340 37324
rect 64647 37284 65340 37312
rect 64647 37281 64659 37284
rect 64601 37275 64659 37281
rect 65334 37272 65340 37284
rect 65392 37272 65398 37324
rect 57517 37247 57575 37253
rect 57517 37213 57529 37247
rect 57563 37213 57575 37247
rect 57517 37207 57575 37213
rect 57701 37247 57759 37253
rect 57701 37213 57713 37247
rect 57747 37244 57759 37247
rect 57790 37244 57796 37256
rect 57747 37216 57796 37244
rect 57747 37213 57759 37216
rect 57701 37207 57759 37213
rect 57532 37176 57560 37207
rect 57790 37204 57796 37216
rect 57848 37244 57854 37256
rect 59998 37244 60004 37256
rect 57848 37216 60004 37244
rect 57848 37204 57854 37216
rect 59998 37204 60004 37216
rect 60056 37204 60062 37256
rect 66898 37204 66904 37256
rect 66956 37244 66962 37256
rect 67085 37247 67143 37253
rect 67085 37244 67097 37247
rect 66956 37216 67097 37244
rect 66956 37204 66962 37216
rect 67085 37213 67097 37216
rect 67131 37213 67143 37247
rect 67085 37207 67143 37213
rect 75362 37204 75368 37256
rect 75420 37204 75426 37256
rect 77297 37247 77355 37253
rect 77297 37213 77309 37247
rect 77343 37213 77355 37247
rect 77297 37207 77355 37213
rect 57974 37176 57980 37188
rect 57532 37148 57980 37176
rect 57974 37136 57980 37148
rect 58032 37136 58038 37188
rect 65978 37176 65984 37188
rect 65826 37148 65984 37176
rect 65978 37136 65984 37148
rect 66036 37136 66042 37188
rect 66916 37176 66944 37204
rect 66088 37148 66944 37176
rect 75273 37179 75331 37185
rect 56778 37068 56784 37120
rect 56836 37108 56842 37120
rect 57330 37108 57336 37120
rect 56836 37080 57336 37108
rect 56836 37068 56842 37080
rect 57330 37068 57336 37080
rect 57388 37108 57394 37120
rect 66088 37117 66116 37148
rect 75273 37145 75285 37179
rect 75319 37176 75331 37179
rect 76098 37176 76104 37188
rect 75319 37148 76104 37176
rect 75319 37145 75331 37148
rect 75273 37139 75331 37145
rect 76098 37136 76104 37148
rect 76156 37176 76162 37188
rect 77312 37176 77340 37207
rect 76156 37148 77340 37176
rect 76156 37136 76162 37148
rect 57609 37111 57667 37117
rect 57609 37108 57621 37111
rect 57388 37080 57621 37108
rect 57388 37068 57394 37080
rect 57609 37077 57621 37080
rect 57655 37077 57667 37111
rect 57609 37071 57667 37077
rect 66073 37111 66131 37117
rect 66073 37077 66085 37111
rect 66119 37077 66131 37111
rect 66073 37071 66131 37077
rect 66530 37068 66536 37120
rect 66588 37068 66594 37120
rect 77478 37068 77484 37120
rect 77536 37068 77542 37120
rect 2024 37018 77924 37040
rect 2024 36966 5794 37018
rect 5846 36966 5858 37018
rect 5910 36966 5922 37018
rect 5974 36966 5986 37018
rect 6038 36966 6050 37018
rect 6102 36966 36514 37018
rect 36566 36966 36578 37018
rect 36630 36966 36642 37018
rect 36694 36966 36706 37018
rect 36758 36966 36770 37018
rect 36822 36966 67234 37018
rect 67286 36966 67298 37018
rect 67350 36966 67362 37018
rect 67414 36966 67426 37018
rect 67478 36966 67490 37018
rect 67542 36966 77924 37018
rect 2024 36944 77924 36966
rect 65334 36864 65340 36916
rect 65392 36904 65398 36916
rect 65429 36907 65487 36913
rect 65429 36904 65441 36907
rect 65392 36876 65441 36904
rect 65392 36864 65398 36876
rect 65429 36873 65441 36876
rect 65475 36873 65487 36907
rect 65429 36867 65487 36873
rect 65978 36864 65984 36916
rect 66036 36904 66042 36916
rect 66073 36907 66131 36913
rect 66073 36904 66085 36907
rect 66036 36876 66085 36904
rect 66036 36864 66042 36876
rect 66073 36873 66085 36876
rect 66119 36873 66131 36907
rect 66073 36867 66131 36873
rect 59998 36796 60004 36848
rect 60056 36796 60062 36848
rect 60366 36796 60372 36848
rect 60424 36796 60430 36848
rect 60737 36839 60795 36845
rect 60737 36805 60749 36839
rect 60783 36836 60795 36839
rect 60918 36836 60924 36848
rect 60783 36808 60924 36836
rect 60783 36805 60795 36808
rect 60737 36799 60795 36805
rect 60918 36796 60924 36808
rect 60976 36796 60982 36848
rect 66530 36836 66536 36848
rect 65904 36808 66536 36836
rect 57974 36728 57980 36780
rect 58032 36768 58038 36780
rect 60182 36768 60188 36780
rect 58032 36740 60188 36768
rect 58032 36728 58038 36740
rect 60182 36728 60188 36740
rect 60240 36728 60246 36780
rect 60274 36728 60280 36780
rect 60332 36728 60338 36780
rect 65610 36728 65616 36780
rect 65668 36728 65674 36780
rect 65794 36728 65800 36780
rect 65852 36728 65858 36780
rect 65904 36777 65932 36808
rect 66530 36796 66536 36808
rect 66588 36796 66594 36848
rect 65889 36771 65947 36777
rect 65889 36737 65901 36771
rect 65935 36737 65947 36771
rect 65889 36731 65947 36737
rect 66162 36728 66168 36780
rect 66220 36768 66226 36780
rect 66990 36768 66996 36780
rect 66220 36740 66996 36768
rect 66220 36728 66226 36740
rect 66990 36728 66996 36740
rect 67048 36728 67054 36780
rect 2024 36474 77924 36496
rect 2024 36422 5134 36474
rect 5186 36422 5198 36474
rect 5250 36422 5262 36474
rect 5314 36422 5326 36474
rect 5378 36422 5390 36474
rect 5442 36422 35854 36474
rect 35906 36422 35918 36474
rect 35970 36422 35982 36474
rect 36034 36422 36046 36474
rect 36098 36422 36110 36474
rect 36162 36422 66574 36474
rect 66626 36422 66638 36474
rect 66690 36422 66702 36474
rect 66754 36422 66766 36474
rect 66818 36422 66830 36474
rect 66882 36422 77924 36474
rect 2024 36400 77924 36422
rect 65610 36320 65616 36372
rect 65668 36360 65674 36372
rect 65978 36360 65984 36372
rect 65668 36332 65984 36360
rect 65668 36320 65674 36332
rect 65978 36320 65984 36332
rect 66036 36360 66042 36372
rect 66625 36363 66683 36369
rect 66625 36360 66637 36363
rect 66036 36332 66637 36360
rect 66036 36320 66042 36332
rect 66625 36329 66637 36332
rect 66671 36329 66683 36363
rect 66625 36323 66683 36329
rect 76466 36320 76472 36372
rect 76524 36320 76530 36372
rect 59998 36252 60004 36304
rect 60056 36252 60062 36304
rect 60461 36295 60519 36301
rect 60461 36261 60473 36295
rect 60507 36292 60519 36295
rect 60645 36295 60703 36301
rect 60645 36292 60657 36295
rect 60507 36264 60657 36292
rect 60507 36261 60519 36264
rect 60461 36255 60519 36261
rect 60645 36261 60657 36264
rect 60691 36261 60703 36295
rect 60645 36255 60703 36261
rect 70765 36295 70823 36301
rect 70765 36261 70777 36295
rect 70811 36261 70823 36295
rect 70765 36255 70823 36261
rect 60016 36224 60044 36252
rect 60093 36227 60151 36233
rect 60093 36224 60105 36227
rect 60016 36196 60105 36224
rect 60093 36193 60105 36196
rect 60139 36193 60151 36227
rect 60093 36187 60151 36193
rect 60182 36184 60188 36236
rect 60240 36184 60246 36236
rect 60274 36184 60280 36236
rect 60332 36184 60338 36236
rect 60918 36184 60924 36236
rect 60976 36224 60982 36236
rect 61013 36227 61071 36233
rect 61013 36224 61025 36227
rect 60976 36196 61025 36224
rect 60976 36184 60982 36196
rect 61013 36193 61025 36196
rect 61059 36224 61071 36227
rect 70780 36224 70808 36255
rect 71682 36224 71688 36236
rect 61059 36196 64874 36224
rect 61059 36193 61071 36196
rect 61013 36187 61071 36193
rect 60001 36159 60059 36165
rect 60001 36125 60013 36159
rect 60047 36125 60059 36159
rect 64846 36156 64874 36196
rect 66548 36196 70624 36224
rect 70780 36196 71688 36224
rect 66548 36165 66576 36196
rect 66533 36159 66591 36165
rect 66533 36156 66545 36159
rect 64846 36128 66545 36156
rect 60001 36119 60059 36125
rect 66533 36125 66545 36128
rect 66579 36125 66591 36159
rect 66533 36119 66591 36125
rect 66717 36159 66775 36165
rect 66717 36125 66729 36159
rect 66763 36156 66775 36159
rect 67082 36156 67088 36168
rect 66763 36128 67088 36156
rect 66763 36125 66775 36128
rect 66717 36119 66775 36125
rect 60016 36088 60044 36119
rect 67082 36116 67088 36128
rect 67140 36116 67146 36168
rect 70596 36165 70624 36196
rect 71682 36184 71688 36196
rect 71740 36224 71746 36236
rect 72697 36227 72755 36233
rect 72697 36224 72709 36227
rect 71740 36196 72709 36224
rect 71740 36184 71746 36196
rect 72697 36193 72709 36196
rect 72743 36193 72755 36227
rect 76374 36224 76380 36236
rect 72697 36187 72755 36193
rect 76208 36196 76380 36224
rect 76208 36168 76236 36196
rect 76374 36184 76380 36196
rect 76432 36184 76438 36236
rect 70581 36159 70639 36165
rect 70581 36125 70593 36159
rect 70627 36156 70639 36159
rect 70627 36128 70808 36156
rect 70627 36125 70639 36128
rect 70581 36119 70639 36125
rect 60366 36088 60372 36100
rect 60016 36060 60372 36088
rect 60366 36048 60372 36060
rect 60424 36088 60430 36100
rect 67100 36088 67128 36116
rect 70670 36088 70676 36100
rect 60424 36060 60688 36088
rect 67100 36060 70676 36088
rect 60424 36048 60430 36060
rect 60550 35980 60556 36032
rect 60608 35980 60614 36032
rect 60660 36020 60688 36060
rect 70670 36048 70676 36060
rect 70728 36048 70734 36100
rect 70780 36088 70808 36128
rect 70854 36116 70860 36168
rect 70912 36156 70918 36168
rect 71038 36156 71044 36168
rect 70912 36128 71044 36156
rect 70912 36116 70918 36128
rect 71038 36116 71044 36128
rect 71096 36116 71102 36168
rect 72789 36159 72847 36165
rect 72789 36125 72801 36159
rect 72835 36156 72847 36159
rect 73154 36156 73160 36168
rect 72835 36128 73160 36156
rect 72835 36125 72847 36128
rect 72789 36119 72847 36125
rect 73154 36116 73160 36128
rect 73212 36116 73218 36168
rect 74074 36116 74080 36168
rect 74132 36116 74138 36168
rect 76190 36116 76196 36168
rect 76248 36116 76254 36168
rect 76282 36116 76288 36168
rect 76340 36116 76346 36168
rect 71130 36088 71136 36100
rect 70780 36060 71136 36088
rect 71130 36048 71136 36060
rect 71188 36048 71194 36100
rect 74353 36091 74411 36097
rect 74353 36057 74365 36091
rect 74399 36057 74411 36091
rect 76101 36091 76159 36097
rect 76101 36088 76113 36091
rect 75578 36060 76113 36088
rect 74353 36051 74411 36057
rect 76101 36057 76113 36060
rect 76147 36057 76159 36091
rect 76101 36051 76159 36057
rect 62114 36020 62120 36032
rect 60660 35992 62120 36020
rect 62114 35980 62120 35992
rect 62172 35980 62178 36032
rect 73157 36023 73215 36029
rect 73157 35989 73169 36023
rect 73203 36020 73215 36023
rect 74368 36020 74396 36051
rect 73203 35992 74396 36020
rect 73203 35989 73215 35992
rect 73157 35983 73215 35989
rect 75822 35980 75828 36032
rect 75880 35980 75886 36032
rect 2024 35930 77924 35952
rect 2024 35878 5794 35930
rect 5846 35878 5858 35930
rect 5910 35878 5922 35930
rect 5974 35878 5986 35930
rect 6038 35878 6050 35930
rect 6102 35878 36514 35930
rect 36566 35878 36578 35930
rect 36630 35878 36642 35930
rect 36694 35878 36706 35930
rect 36758 35878 36770 35930
rect 36822 35878 67234 35930
rect 67286 35878 67298 35930
rect 67350 35878 67362 35930
rect 67414 35878 67426 35930
rect 67478 35878 67490 35930
rect 67542 35878 77924 35930
rect 2024 35856 77924 35878
rect 63494 35816 63500 35828
rect 60384 35788 63500 35816
rect 56689 35683 56747 35689
rect 56689 35649 56701 35683
rect 56735 35680 56747 35683
rect 57425 35683 57483 35689
rect 57425 35680 57437 35683
rect 56735 35652 57437 35680
rect 56735 35649 56747 35652
rect 56689 35643 56747 35649
rect 57425 35649 57437 35652
rect 57471 35649 57483 35683
rect 57425 35643 57483 35649
rect 58066 35640 58072 35692
rect 58124 35680 58130 35692
rect 60274 35680 60280 35692
rect 58124 35652 60280 35680
rect 58124 35640 58130 35652
rect 60274 35640 60280 35652
rect 60332 35640 60338 35692
rect 60384 35624 60412 35788
rect 63494 35776 63500 35788
rect 63552 35776 63558 35828
rect 73154 35776 73160 35828
rect 73212 35816 73218 35828
rect 74353 35819 74411 35825
rect 74353 35816 74365 35819
rect 73212 35788 74365 35816
rect 73212 35776 73218 35788
rect 74353 35785 74365 35788
rect 74399 35785 74411 35819
rect 74353 35779 74411 35785
rect 60550 35708 60556 35760
rect 60608 35748 60614 35760
rect 60645 35751 60703 35757
rect 60645 35748 60657 35751
rect 60608 35720 60657 35748
rect 60608 35708 60614 35720
rect 60645 35717 60657 35720
rect 60691 35717 60703 35751
rect 62301 35751 62359 35757
rect 62301 35748 62313 35751
rect 61870 35720 62313 35748
rect 60645 35711 60703 35717
rect 62301 35717 62313 35720
rect 62347 35717 62359 35751
rect 62301 35711 62359 35717
rect 70670 35708 70676 35760
rect 70728 35748 70734 35760
rect 70728 35720 71268 35748
rect 70728 35708 70734 35720
rect 62393 35683 62451 35689
rect 62393 35680 62405 35683
rect 61856 35652 62405 35680
rect 56778 35572 56784 35624
rect 56836 35572 56842 35624
rect 60366 35572 60372 35624
rect 60424 35572 60430 35624
rect 61856 35612 61884 35652
rect 62393 35649 62405 35652
rect 62439 35680 62451 35683
rect 66162 35680 66168 35692
rect 62439 35652 66168 35680
rect 62439 35649 62451 35652
rect 62393 35643 62451 35649
rect 66162 35640 66168 35652
rect 66220 35640 66226 35692
rect 71130 35640 71136 35692
rect 71188 35640 71194 35692
rect 71240 35689 71268 35720
rect 71225 35683 71283 35689
rect 71225 35649 71237 35683
rect 71271 35649 71283 35683
rect 71225 35643 71283 35649
rect 71682 35640 71688 35692
rect 71740 35640 71746 35692
rect 74997 35683 75055 35689
rect 74997 35649 75009 35683
rect 75043 35680 75055 35683
rect 75822 35680 75828 35692
rect 75043 35652 75828 35680
rect 75043 35649 75055 35652
rect 74997 35643 75055 35649
rect 75822 35640 75828 35652
rect 75880 35640 75886 35692
rect 60476 35584 61884 35612
rect 58342 35504 58348 35556
rect 58400 35544 58406 35556
rect 60476 35544 60504 35584
rect 62114 35572 62120 35624
rect 62172 35572 62178 35624
rect 70118 35572 70124 35624
rect 70176 35572 70182 35624
rect 70765 35615 70823 35621
rect 70765 35581 70777 35615
rect 70811 35612 70823 35615
rect 70949 35615 71007 35621
rect 70949 35612 70961 35615
rect 70811 35584 70961 35612
rect 70811 35581 70823 35584
rect 70765 35575 70823 35581
rect 70949 35581 70961 35584
rect 70995 35581 71007 35615
rect 70949 35575 71007 35581
rect 71041 35615 71099 35621
rect 71041 35581 71053 35615
rect 71087 35581 71099 35615
rect 71041 35575 71099 35581
rect 71409 35615 71467 35621
rect 71409 35581 71421 35615
rect 71455 35612 71467 35615
rect 71869 35615 71927 35621
rect 71869 35612 71881 35615
rect 71455 35584 71881 35612
rect 71455 35581 71467 35584
rect 71409 35575 71467 35581
rect 71869 35581 71881 35584
rect 71915 35581 71927 35615
rect 71869 35575 71927 35581
rect 58400 35516 60504 35544
rect 58400 35504 58406 35516
rect 70670 35504 70676 35556
rect 70728 35544 70734 35556
rect 71056 35544 71084 35575
rect 70728 35516 71084 35544
rect 70728 35504 70734 35516
rect 1210 35436 1216 35488
rect 1268 35476 1274 35488
rect 2317 35479 2375 35485
rect 2317 35476 2329 35479
rect 1268 35448 2329 35476
rect 1268 35436 1274 35448
rect 2317 35445 2329 35448
rect 2363 35445 2375 35479
rect 2317 35439 2375 35445
rect 56410 35436 56416 35488
rect 56468 35436 56474 35488
rect 71314 35436 71320 35488
rect 71372 35476 71378 35488
rect 71501 35479 71559 35485
rect 71501 35476 71513 35479
rect 71372 35448 71513 35476
rect 71372 35436 71378 35448
rect 71501 35445 71513 35448
rect 71547 35445 71559 35479
rect 71501 35439 71559 35445
rect 2024 35386 77924 35408
rect 2024 35334 5134 35386
rect 5186 35334 5198 35386
rect 5250 35334 5262 35386
rect 5314 35334 5326 35386
rect 5378 35334 5390 35386
rect 5442 35334 35854 35386
rect 35906 35334 35918 35386
rect 35970 35334 35982 35386
rect 36034 35334 36046 35386
rect 36098 35334 36110 35386
rect 36162 35334 66574 35386
rect 66626 35334 66638 35386
rect 66690 35334 66702 35386
rect 66754 35334 66766 35386
rect 66818 35334 66830 35386
rect 66882 35334 77924 35386
rect 2024 35312 77924 35334
rect 56410 35232 56416 35284
rect 56468 35272 56474 35284
rect 56578 35275 56636 35281
rect 56578 35272 56590 35275
rect 56468 35244 56590 35272
rect 56468 35232 56474 35244
rect 56578 35241 56590 35244
rect 56624 35241 56636 35275
rect 56578 35235 56636 35241
rect 58066 35232 58072 35284
rect 58124 35232 58130 35284
rect 70854 35232 70860 35284
rect 70912 35272 70918 35284
rect 70949 35275 71007 35281
rect 70949 35272 70961 35275
rect 70912 35244 70961 35272
rect 70912 35232 70918 35244
rect 70949 35241 70961 35244
rect 70995 35241 71007 35275
rect 70949 35235 71007 35241
rect 56321 35139 56379 35145
rect 56321 35105 56333 35139
rect 56367 35136 56379 35139
rect 60366 35136 60372 35148
rect 56367 35108 60372 35136
rect 56367 35105 56379 35108
rect 56321 35099 56379 35105
rect 60366 35096 60372 35108
rect 60424 35096 60430 35148
rect 70118 35096 70124 35148
rect 70176 35136 70182 35148
rect 70176 35108 70808 35136
rect 70176 35096 70182 35108
rect 58342 35028 58348 35080
rect 58400 35028 58406 35080
rect 66990 35028 66996 35080
rect 67048 35068 67054 35080
rect 70670 35068 70676 35080
rect 67048 35040 70676 35068
rect 67048 35028 67054 35040
rect 70670 35028 70676 35040
rect 70728 35028 70734 35080
rect 70780 35077 70808 35108
rect 70765 35071 70823 35077
rect 70765 35037 70777 35071
rect 70811 35037 70823 35071
rect 70765 35031 70823 35037
rect 58253 35003 58311 35009
rect 58253 35000 58265 35003
rect 57822 34972 58265 35000
rect 58253 34969 58265 34972
rect 58299 34969 58311 35003
rect 58253 34963 58311 34969
rect 2024 34842 77924 34864
rect 2024 34790 5794 34842
rect 5846 34790 5858 34842
rect 5910 34790 5922 34842
rect 5974 34790 5986 34842
rect 6038 34790 6050 34842
rect 6102 34790 36514 34842
rect 36566 34790 36578 34842
rect 36630 34790 36642 34842
rect 36694 34790 36706 34842
rect 36758 34790 36770 34842
rect 36822 34790 67234 34842
rect 67286 34790 67298 34842
rect 67350 34790 67362 34842
rect 67414 34790 67426 34842
rect 67478 34790 67490 34842
rect 67542 34790 77924 34842
rect 2024 34768 77924 34790
rect 68922 34688 68928 34740
rect 68980 34728 68986 34740
rect 68980 34700 71636 34728
rect 68980 34688 68986 34700
rect 70302 34620 70308 34672
rect 70360 34620 70366 34672
rect 71314 34620 71320 34672
rect 71372 34620 71378 34672
rect 71608 34660 71636 34700
rect 74074 34660 74080 34672
rect 71608 34632 74080 34660
rect 65889 34595 65947 34601
rect 65889 34561 65901 34595
rect 65935 34592 65947 34595
rect 66349 34595 66407 34601
rect 66349 34592 66361 34595
rect 65935 34564 66361 34592
rect 65935 34561 65947 34564
rect 65889 34555 65947 34561
rect 66349 34561 66361 34564
rect 66395 34561 66407 34595
rect 66349 34555 66407 34561
rect 66990 34552 66996 34604
rect 67048 34552 67054 34604
rect 71608 34601 71636 34632
rect 74074 34620 74080 34632
rect 74132 34620 74138 34672
rect 76190 34660 76196 34672
rect 74506 34632 76196 34660
rect 71593 34595 71651 34601
rect 71593 34561 71605 34595
rect 71639 34561 71651 34595
rect 71593 34555 71651 34561
rect 72145 34595 72203 34601
rect 72145 34561 72157 34595
rect 72191 34592 72203 34595
rect 74506 34592 74534 34632
rect 76190 34620 76196 34632
rect 76248 34660 76254 34672
rect 77297 34663 77355 34669
rect 77297 34660 77309 34663
rect 76248 34632 77309 34660
rect 76248 34620 76254 34632
rect 77297 34629 77309 34632
rect 77343 34629 77355 34663
rect 77297 34623 77355 34629
rect 72191 34564 74534 34592
rect 72191 34561 72203 34564
rect 72145 34555 72203 34561
rect 77478 34552 77484 34604
rect 77536 34552 77542 34604
rect 65978 34484 65984 34536
rect 66036 34484 66042 34536
rect 69845 34527 69903 34533
rect 69845 34493 69857 34527
rect 69891 34524 69903 34527
rect 70118 34524 70124 34536
rect 69891 34496 70124 34524
rect 69891 34493 69903 34496
rect 69845 34487 69903 34493
rect 70118 34484 70124 34496
rect 70176 34484 70182 34536
rect 71866 34484 71872 34536
rect 71924 34484 71930 34536
rect 66165 34391 66223 34397
rect 66165 34357 66177 34391
rect 66211 34388 66223 34391
rect 68002 34388 68008 34400
rect 66211 34360 68008 34388
rect 66211 34357 66223 34360
rect 66165 34351 66223 34357
rect 68002 34348 68008 34360
rect 68060 34348 68066 34400
rect 2024 34298 77924 34320
rect 2024 34246 5134 34298
rect 5186 34246 5198 34298
rect 5250 34246 5262 34298
rect 5314 34246 5326 34298
rect 5378 34246 5390 34298
rect 5442 34246 35854 34298
rect 35906 34246 35918 34298
rect 35970 34246 35982 34298
rect 36034 34246 36046 34298
rect 36098 34246 36110 34298
rect 36162 34246 66574 34298
rect 66626 34246 66638 34298
rect 66690 34246 66702 34298
rect 66754 34246 66766 34298
rect 66818 34246 66830 34298
rect 66882 34246 77924 34298
rect 2024 34224 77924 34246
rect 66533 34187 66591 34193
rect 66533 34153 66545 34187
rect 66579 34184 66591 34187
rect 66990 34184 66996 34196
rect 66579 34156 66996 34184
rect 66579 34153 66591 34156
rect 66533 34147 66591 34153
rect 66990 34144 66996 34156
rect 67048 34144 67054 34196
rect 70302 34144 70308 34196
rect 70360 34184 70366 34196
rect 70949 34187 71007 34193
rect 70949 34184 70961 34187
rect 70360 34156 70961 34184
rect 70360 34144 70366 34156
rect 70949 34153 70961 34156
rect 70995 34153 71007 34187
rect 70949 34147 71007 34153
rect 68002 34008 68008 34060
rect 68060 34008 68066 34060
rect 68281 34051 68339 34057
rect 68281 34017 68293 34051
rect 68327 34048 68339 34051
rect 68922 34048 68928 34060
rect 68327 34020 68928 34048
rect 68327 34017 68339 34020
rect 68281 34011 68339 34017
rect 68922 34008 68928 34020
rect 68980 34008 68986 34060
rect 66898 33940 66904 33992
rect 66956 33940 66962 33992
rect 71041 33983 71099 33989
rect 71041 33949 71053 33983
rect 71087 33980 71099 33983
rect 71866 33980 71872 33992
rect 71087 33952 71872 33980
rect 71087 33949 71099 33952
rect 71041 33943 71099 33949
rect 66254 33804 66260 33856
rect 66312 33844 66318 33856
rect 71056 33844 71084 33943
rect 71866 33940 71872 33952
rect 71924 33940 71930 33992
rect 66312 33816 71084 33844
rect 66312 33804 66318 33816
rect 2024 33754 77924 33776
rect 2024 33702 5794 33754
rect 5846 33702 5858 33754
rect 5910 33702 5922 33754
rect 5974 33702 5986 33754
rect 6038 33702 6050 33754
rect 6102 33702 36514 33754
rect 36566 33702 36578 33754
rect 36630 33702 36642 33754
rect 36694 33702 36706 33754
rect 36758 33702 36770 33754
rect 36822 33702 67234 33754
rect 67286 33702 67298 33754
rect 67350 33702 67362 33754
rect 67414 33702 67426 33754
rect 67478 33702 67490 33754
rect 67542 33702 77924 33754
rect 2024 33680 77924 33702
rect 66898 33600 66904 33652
rect 66956 33600 66962 33652
rect 66254 33464 66260 33516
rect 66312 33504 66318 33516
rect 66809 33507 66867 33513
rect 66809 33504 66821 33507
rect 66312 33476 66821 33504
rect 66312 33464 66318 33476
rect 66809 33473 66821 33476
rect 66855 33473 66867 33507
rect 66809 33467 66867 33473
rect 2024 33210 77924 33232
rect 2024 33158 5134 33210
rect 5186 33158 5198 33210
rect 5250 33158 5262 33210
rect 5314 33158 5326 33210
rect 5378 33158 5390 33210
rect 5442 33158 35854 33210
rect 35906 33158 35918 33210
rect 35970 33158 35982 33210
rect 36034 33158 36046 33210
rect 36098 33158 36110 33210
rect 36162 33158 66574 33210
rect 66626 33158 66638 33210
rect 66690 33158 66702 33210
rect 66754 33158 66766 33210
rect 66818 33158 66830 33210
rect 66882 33158 77924 33210
rect 2024 33136 77924 33158
rect 2024 32666 77924 32688
rect 2024 32614 5794 32666
rect 5846 32614 5858 32666
rect 5910 32614 5922 32666
rect 5974 32614 5986 32666
rect 6038 32614 6050 32666
rect 6102 32614 36514 32666
rect 36566 32614 36578 32666
rect 36630 32614 36642 32666
rect 36694 32614 36706 32666
rect 36758 32614 36770 32666
rect 36822 32614 67234 32666
rect 67286 32614 67298 32666
rect 67350 32614 67362 32666
rect 67414 32614 67426 32666
rect 67478 32614 67490 32666
rect 67542 32614 77924 32666
rect 2024 32592 77924 32614
rect 1210 32172 1216 32224
rect 1268 32212 1274 32224
rect 2317 32215 2375 32221
rect 2317 32212 2329 32215
rect 1268 32184 2329 32212
rect 1268 32172 1274 32184
rect 2317 32181 2329 32184
rect 2363 32181 2375 32215
rect 2317 32175 2375 32181
rect 2024 32122 77924 32144
rect 2024 32070 5134 32122
rect 5186 32070 5198 32122
rect 5250 32070 5262 32122
rect 5314 32070 5326 32122
rect 5378 32070 5390 32122
rect 5442 32070 35854 32122
rect 35906 32070 35918 32122
rect 35970 32070 35982 32122
rect 36034 32070 36046 32122
rect 36098 32070 36110 32122
rect 36162 32070 66574 32122
rect 66626 32070 66638 32122
rect 66690 32070 66702 32122
rect 66754 32070 66766 32122
rect 66818 32070 66830 32122
rect 66882 32070 77924 32122
rect 2024 32048 77924 32070
rect 2024 31578 77924 31600
rect 2024 31526 5794 31578
rect 5846 31526 5858 31578
rect 5910 31526 5922 31578
rect 5974 31526 5986 31578
rect 6038 31526 6050 31578
rect 6102 31526 36514 31578
rect 36566 31526 36578 31578
rect 36630 31526 36642 31578
rect 36694 31526 36706 31578
rect 36758 31526 36770 31578
rect 36822 31526 67234 31578
rect 67286 31526 67298 31578
rect 67350 31526 67362 31578
rect 67414 31526 67426 31578
rect 67478 31526 67490 31578
rect 67542 31526 77924 31578
rect 2024 31504 77924 31526
rect 2024 31034 77924 31056
rect 2024 30982 5134 31034
rect 5186 30982 5198 31034
rect 5250 30982 5262 31034
rect 5314 30982 5326 31034
rect 5378 30982 5390 31034
rect 5442 30982 35854 31034
rect 35906 30982 35918 31034
rect 35970 30982 35982 31034
rect 36034 30982 36046 31034
rect 36098 30982 36110 31034
rect 36162 30982 66574 31034
rect 66626 30982 66638 31034
rect 66690 30982 66702 31034
rect 66754 30982 66766 31034
rect 66818 30982 66830 31034
rect 66882 30982 77924 31034
rect 2024 30960 77924 30982
rect 2024 30490 77924 30512
rect 2024 30438 5794 30490
rect 5846 30438 5858 30490
rect 5910 30438 5922 30490
rect 5974 30438 5986 30490
rect 6038 30438 6050 30490
rect 6102 30438 36514 30490
rect 36566 30438 36578 30490
rect 36630 30438 36642 30490
rect 36694 30438 36706 30490
rect 36758 30438 36770 30490
rect 36822 30438 67234 30490
rect 67286 30438 67298 30490
rect 67350 30438 67362 30490
rect 67414 30438 67426 30490
rect 67478 30438 67490 30490
rect 67542 30438 77924 30490
rect 2024 30416 77924 30438
rect 2024 29946 77924 29968
rect 2024 29894 5134 29946
rect 5186 29894 5198 29946
rect 5250 29894 5262 29946
rect 5314 29894 5326 29946
rect 5378 29894 5390 29946
rect 5442 29894 35854 29946
rect 35906 29894 35918 29946
rect 35970 29894 35982 29946
rect 36034 29894 36046 29946
rect 36098 29894 36110 29946
rect 36162 29894 66574 29946
rect 66626 29894 66638 29946
rect 66690 29894 66702 29946
rect 66754 29894 66766 29946
rect 66818 29894 66830 29946
rect 66882 29894 77924 29946
rect 2024 29872 77924 29894
rect 2024 29402 77924 29424
rect 2024 29350 5794 29402
rect 5846 29350 5858 29402
rect 5910 29350 5922 29402
rect 5974 29350 5986 29402
rect 6038 29350 6050 29402
rect 6102 29350 36514 29402
rect 36566 29350 36578 29402
rect 36630 29350 36642 29402
rect 36694 29350 36706 29402
rect 36758 29350 36770 29402
rect 36822 29350 67234 29402
rect 67286 29350 67298 29402
rect 67350 29350 67362 29402
rect 67414 29350 67426 29402
rect 67478 29350 67490 29402
rect 67542 29350 77924 29402
rect 2024 29328 77924 29350
rect 2314 28976 2320 29028
rect 2372 28976 2378 29028
rect 2024 28858 77924 28880
rect 2024 28806 5134 28858
rect 5186 28806 5198 28858
rect 5250 28806 5262 28858
rect 5314 28806 5326 28858
rect 5378 28806 5390 28858
rect 5442 28806 35854 28858
rect 35906 28806 35918 28858
rect 35970 28806 35982 28858
rect 36034 28806 36046 28858
rect 36098 28806 36110 28858
rect 36162 28806 66574 28858
rect 66626 28806 66638 28858
rect 66690 28806 66702 28858
rect 66754 28806 66766 28858
rect 66818 28806 66830 28858
rect 66882 28806 77924 28858
rect 2024 28784 77924 28806
rect 2024 28314 77924 28336
rect 2024 28262 5794 28314
rect 5846 28262 5858 28314
rect 5910 28262 5922 28314
rect 5974 28262 5986 28314
rect 6038 28262 6050 28314
rect 6102 28262 36514 28314
rect 36566 28262 36578 28314
rect 36630 28262 36642 28314
rect 36694 28262 36706 28314
rect 36758 28262 36770 28314
rect 36822 28262 67234 28314
rect 67286 28262 67298 28314
rect 67350 28262 67362 28314
rect 67414 28262 67426 28314
rect 67478 28262 67490 28314
rect 67542 28262 77924 28314
rect 2024 28240 77924 28262
rect 1210 27956 1216 28008
rect 1268 27996 1274 28008
rect 2317 27999 2375 28005
rect 2317 27996 2329 27999
rect 1268 27968 2329 27996
rect 1268 27956 1274 27968
rect 2317 27965 2329 27968
rect 2363 27965 2375 27999
rect 2317 27959 2375 27965
rect 2024 27770 77924 27792
rect 2024 27718 5134 27770
rect 5186 27718 5198 27770
rect 5250 27718 5262 27770
rect 5314 27718 5326 27770
rect 5378 27718 5390 27770
rect 5442 27718 35854 27770
rect 35906 27718 35918 27770
rect 35970 27718 35982 27770
rect 36034 27718 36046 27770
rect 36098 27718 36110 27770
rect 36162 27718 66574 27770
rect 66626 27718 66638 27770
rect 66690 27718 66702 27770
rect 66754 27718 66766 27770
rect 66818 27718 66830 27770
rect 66882 27718 77924 27770
rect 2024 27696 77924 27718
rect 2024 27226 77924 27248
rect 2024 27174 5794 27226
rect 5846 27174 5858 27226
rect 5910 27174 5922 27226
rect 5974 27174 5986 27226
rect 6038 27174 6050 27226
rect 6102 27174 36514 27226
rect 36566 27174 36578 27226
rect 36630 27174 36642 27226
rect 36694 27174 36706 27226
rect 36758 27174 36770 27226
rect 36822 27174 67234 27226
rect 67286 27174 67298 27226
rect 67350 27174 67362 27226
rect 67414 27174 67426 27226
rect 67478 27174 67490 27226
rect 67542 27174 77924 27226
rect 2024 27152 77924 27174
rect 1210 26732 1216 26784
rect 1268 26772 1274 26784
rect 2317 26775 2375 26781
rect 2317 26772 2329 26775
rect 1268 26744 2329 26772
rect 1268 26732 1274 26744
rect 2317 26741 2329 26744
rect 2363 26741 2375 26775
rect 2317 26735 2375 26741
rect 2024 26682 77924 26704
rect 2024 26630 5134 26682
rect 5186 26630 5198 26682
rect 5250 26630 5262 26682
rect 5314 26630 5326 26682
rect 5378 26630 5390 26682
rect 5442 26630 35854 26682
rect 35906 26630 35918 26682
rect 35970 26630 35982 26682
rect 36034 26630 36046 26682
rect 36098 26630 36110 26682
rect 36162 26630 66574 26682
rect 66626 26630 66638 26682
rect 66690 26630 66702 26682
rect 66754 26630 66766 26682
rect 66818 26630 66830 26682
rect 66882 26630 77924 26682
rect 2024 26608 77924 26630
rect 2314 26324 2320 26376
rect 2372 26324 2378 26376
rect 2024 26138 77924 26160
rect 2024 26086 5794 26138
rect 5846 26086 5858 26138
rect 5910 26086 5922 26138
rect 5974 26086 5986 26138
rect 6038 26086 6050 26138
rect 6102 26086 36514 26138
rect 36566 26086 36578 26138
rect 36630 26086 36642 26138
rect 36694 26086 36706 26138
rect 36758 26086 36770 26138
rect 36822 26086 67234 26138
rect 67286 26086 67298 26138
rect 67350 26086 67362 26138
rect 67414 26086 67426 26138
rect 67478 26086 67490 26138
rect 67542 26086 77924 26138
rect 2024 26064 77924 26086
rect 2024 25594 77924 25616
rect 2024 25542 5134 25594
rect 5186 25542 5198 25594
rect 5250 25542 5262 25594
rect 5314 25542 5326 25594
rect 5378 25542 5390 25594
rect 5442 25542 35854 25594
rect 35906 25542 35918 25594
rect 35970 25542 35982 25594
rect 36034 25542 36046 25594
rect 36098 25542 36110 25594
rect 36162 25542 66574 25594
rect 66626 25542 66638 25594
rect 66690 25542 66702 25594
rect 66754 25542 66766 25594
rect 66818 25542 66830 25594
rect 66882 25542 77924 25594
rect 2024 25520 77924 25542
rect 2024 25050 77924 25072
rect 2024 24998 5794 25050
rect 5846 24998 5858 25050
rect 5910 24998 5922 25050
rect 5974 24998 5986 25050
rect 6038 24998 6050 25050
rect 6102 24998 36514 25050
rect 36566 24998 36578 25050
rect 36630 24998 36642 25050
rect 36694 24998 36706 25050
rect 36758 24998 36770 25050
rect 36822 24998 67234 25050
rect 67286 24998 67298 25050
rect 67350 24998 67362 25050
rect 67414 24998 67426 25050
rect 67478 24998 67490 25050
rect 67542 24998 77924 25050
rect 2024 24976 77924 24998
rect 2024 24506 77924 24528
rect 2024 24454 5134 24506
rect 5186 24454 5198 24506
rect 5250 24454 5262 24506
rect 5314 24454 5326 24506
rect 5378 24454 5390 24506
rect 5442 24454 35854 24506
rect 35906 24454 35918 24506
rect 35970 24454 35982 24506
rect 36034 24454 36046 24506
rect 36098 24454 36110 24506
rect 36162 24454 66574 24506
rect 66626 24454 66638 24506
rect 66690 24454 66702 24506
rect 66754 24454 66766 24506
rect 66818 24454 66830 24506
rect 66882 24454 77924 24506
rect 2024 24432 77924 24454
rect 2024 23962 77924 23984
rect 2024 23910 5794 23962
rect 5846 23910 5858 23962
rect 5910 23910 5922 23962
rect 5974 23910 5986 23962
rect 6038 23910 6050 23962
rect 6102 23910 36514 23962
rect 36566 23910 36578 23962
rect 36630 23910 36642 23962
rect 36694 23910 36706 23962
rect 36758 23910 36770 23962
rect 36822 23910 67234 23962
rect 67286 23910 67298 23962
rect 67350 23910 67362 23962
rect 67414 23910 67426 23962
rect 67478 23910 67490 23962
rect 67542 23910 77924 23962
rect 2024 23888 77924 23910
rect 2314 23468 2320 23520
rect 2372 23468 2378 23520
rect 2024 23418 77924 23440
rect 2024 23366 5134 23418
rect 5186 23366 5198 23418
rect 5250 23366 5262 23418
rect 5314 23366 5326 23418
rect 5378 23366 5390 23418
rect 5442 23366 35854 23418
rect 35906 23366 35918 23418
rect 35970 23366 35982 23418
rect 36034 23366 36046 23418
rect 36098 23366 36110 23418
rect 36162 23366 66574 23418
rect 66626 23366 66638 23418
rect 66690 23366 66702 23418
rect 66754 23366 66766 23418
rect 66818 23366 66830 23418
rect 66882 23366 77924 23418
rect 2024 23344 77924 23366
rect 2024 22874 77924 22896
rect 2024 22822 5794 22874
rect 5846 22822 5858 22874
rect 5910 22822 5922 22874
rect 5974 22822 5986 22874
rect 6038 22822 6050 22874
rect 6102 22822 36514 22874
rect 36566 22822 36578 22874
rect 36630 22822 36642 22874
rect 36694 22822 36706 22874
rect 36758 22822 36770 22874
rect 36822 22822 67234 22874
rect 67286 22822 67298 22874
rect 67350 22822 67362 22874
rect 67414 22822 67426 22874
rect 67478 22822 67490 22874
rect 67542 22822 77924 22874
rect 2024 22800 77924 22822
rect 2024 22330 77924 22352
rect 2024 22278 5134 22330
rect 5186 22278 5198 22330
rect 5250 22278 5262 22330
rect 5314 22278 5326 22330
rect 5378 22278 5390 22330
rect 5442 22278 35854 22330
rect 35906 22278 35918 22330
rect 35970 22278 35982 22330
rect 36034 22278 36046 22330
rect 36098 22278 36110 22330
rect 36162 22278 66574 22330
rect 66626 22278 66638 22330
rect 66690 22278 66702 22330
rect 66754 22278 66766 22330
rect 66818 22278 66830 22330
rect 66882 22278 77924 22330
rect 2024 22256 77924 22278
rect 2024 21786 77924 21808
rect 2024 21734 5794 21786
rect 5846 21734 5858 21786
rect 5910 21734 5922 21786
rect 5974 21734 5986 21786
rect 6038 21734 6050 21786
rect 6102 21734 36514 21786
rect 36566 21734 36578 21786
rect 36630 21734 36642 21786
rect 36694 21734 36706 21786
rect 36758 21734 36770 21786
rect 36822 21734 67234 21786
rect 67286 21734 67298 21786
rect 67350 21734 67362 21786
rect 67414 21734 67426 21786
rect 67478 21734 67490 21786
rect 67542 21734 77924 21786
rect 2024 21712 77924 21734
rect 77570 21292 77576 21344
rect 77628 21292 77634 21344
rect 2024 21242 77924 21264
rect 2024 21190 5134 21242
rect 5186 21190 5198 21242
rect 5250 21190 5262 21242
rect 5314 21190 5326 21242
rect 5378 21190 5390 21242
rect 5442 21190 35854 21242
rect 35906 21190 35918 21242
rect 35970 21190 35982 21242
rect 36034 21190 36046 21242
rect 36098 21190 36110 21242
rect 36162 21190 66574 21242
rect 66626 21190 66638 21242
rect 66690 21190 66702 21242
rect 66754 21190 66766 21242
rect 66818 21190 66830 21242
rect 66882 21190 77924 21242
rect 2024 21168 77924 21190
rect 2024 20698 77924 20720
rect 2024 20646 5794 20698
rect 5846 20646 5858 20698
rect 5910 20646 5922 20698
rect 5974 20646 5986 20698
rect 6038 20646 6050 20698
rect 6102 20646 36514 20698
rect 36566 20646 36578 20698
rect 36630 20646 36642 20698
rect 36694 20646 36706 20698
rect 36758 20646 36770 20698
rect 36822 20646 67234 20698
rect 67286 20646 67298 20698
rect 67350 20646 67362 20698
rect 67414 20646 67426 20698
rect 67478 20646 67490 20698
rect 67542 20646 77924 20698
rect 2024 20624 77924 20646
rect 2024 20154 77924 20176
rect 2024 20102 5134 20154
rect 5186 20102 5198 20154
rect 5250 20102 5262 20154
rect 5314 20102 5326 20154
rect 5378 20102 5390 20154
rect 5442 20102 35854 20154
rect 35906 20102 35918 20154
rect 35970 20102 35982 20154
rect 36034 20102 36046 20154
rect 36098 20102 36110 20154
rect 36162 20102 66574 20154
rect 66626 20102 66638 20154
rect 66690 20102 66702 20154
rect 66754 20102 66766 20154
rect 66818 20102 66830 20154
rect 66882 20102 77924 20154
rect 2024 20080 77924 20102
rect 2024 19610 77924 19632
rect 2024 19558 5794 19610
rect 5846 19558 5858 19610
rect 5910 19558 5922 19610
rect 5974 19558 5986 19610
rect 6038 19558 6050 19610
rect 6102 19558 36514 19610
rect 36566 19558 36578 19610
rect 36630 19558 36642 19610
rect 36694 19558 36706 19610
rect 36758 19558 36770 19610
rect 36822 19558 67234 19610
rect 67286 19558 67298 19610
rect 67350 19558 67362 19610
rect 67414 19558 67426 19610
rect 67478 19558 67490 19610
rect 67542 19558 77924 19610
rect 2024 19536 77924 19558
rect 2024 19066 77924 19088
rect 2024 19014 5134 19066
rect 5186 19014 5198 19066
rect 5250 19014 5262 19066
rect 5314 19014 5326 19066
rect 5378 19014 5390 19066
rect 5442 19014 35854 19066
rect 35906 19014 35918 19066
rect 35970 19014 35982 19066
rect 36034 19014 36046 19066
rect 36098 19014 36110 19066
rect 36162 19014 66574 19066
rect 66626 19014 66638 19066
rect 66690 19014 66702 19066
rect 66754 19014 66766 19066
rect 66818 19014 66830 19066
rect 66882 19014 77924 19066
rect 2024 18992 77924 19014
rect 2024 18522 77924 18544
rect 2024 18470 5794 18522
rect 5846 18470 5858 18522
rect 5910 18470 5922 18522
rect 5974 18470 5986 18522
rect 6038 18470 6050 18522
rect 6102 18470 36514 18522
rect 36566 18470 36578 18522
rect 36630 18470 36642 18522
rect 36694 18470 36706 18522
rect 36758 18470 36770 18522
rect 36822 18470 67234 18522
rect 67286 18470 67298 18522
rect 67350 18470 67362 18522
rect 67414 18470 67426 18522
rect 67478 18470 67490 18522
rect 67542 18470 77924 18522
rect 2024 18448 77924 18470
rect 2024 17978 77924 18000
rect 2024 17926 5134 17978
rect 5186 17926 5198 17978
rect 5250 17926 5262 17978
rect 5314 17926 5326 17978
rect 5378 17926 5390 17978
rect 5442 17926 35854 17978
rect 35906 17926 35918 17978
rect 35970 17926 35982 17978
rect 36034 17926 36046 17978
rect 36098 17926 36110 17978
rect 36162 17926 66574 17978
rect 66626 17926 66638 17978
rect 66690 17926 66702 17978
rect 66754 17926 66766 17978
rect 66818 17926 66830 17978
rect 66882 17926 77924 17978
rect 2024 17904 77924 17926
rect 2024 17434 77924 17456
rect 2024 17382 5794 17434
rect 5846 17382 5858 17434
rect 5910 17382 5922 17434
rect 5974 17382 5986 17434
rect 6038 17382 6050 17434
rect 6102 17382 36514 17434
rect 36566 17382 36578 17434
rect 36630 17382 36642 17434
rect 36694 17382 36706 17434
rect 36758 17382 36770 17434
rect 36822 17382 67234 17434
rect 67286 17382 67298 17434
rect 67350 17382 67362 17434
rect 67414 17382 67426 17434
rect 67478 17382 67490 17434
rect 67542 17382 77924 17434
rect 2024 17360 77924 17382
rect 2024 16890 77924 16912
rect 2024 16838 5134 16890
rect 5186 16838 5198 16890
rect 5250 16838 5262 16890
rect 5314 16838 5326 16890
rect 5378 16838 5390 16890
rect 5442 16838 35854 16890
rect 35906 16838 35918 16890
rect 35970 16838 35982 16890
rect 36034 16838 36046 16890
rect 36098 16838 36110 16890
rect 36162 16838 66574 16890
rect 66626 16838 66638 16890
rect 66690 16838 66702 16890
rect 66754 16838 66766 16890
rect 66818 16838 66830 16890
rect 66882 16838 77924 16890
rect 2024 16816 77924 16838
rect 77570 16600 77576 16652
rect 77628 16600 77634 16652
rect 2024 16346 77924 16368
rect 2024 16294 5794 16346
rect 5846 16294 5858 16346
rect 5910 16294 5922 16346
rect 5974 16294 5986 16346
rect 6038 16294 6050 16346
rect 6102 16294 36514 16346
rect 36566 16294 36578 16346
rect 36630 16294 36642 16346
rect 36694 16294 36706 16346
rect 36758 16294 36770 16346
rect 36822 16294 67234 16346
rect 67286 16294 67298 16346
rect 67350 16294 67362 16346
rect 67414 16294 67426 16346
rect 67478 16294 67490 16346
rect 67542 16294 77924 16346
rect 2024 16272 77924 16294
rect 2024 15802 77924 15824
rect 2024 15750 5134 15802
rect 5186 15750 5198 15802
rect 5250 15750 5262 15802
rect 5314 15750 5326 15802
rect 5378 15750 5390 15802
rect 5442 15750 35854 15802
rect 35906 15750 35918 15802
rect 35970 15750 35982 15802
rect 36034 15750 36046 15802
rect 36098 15750 36110 15802
rect 36162 15750 66574 15802
rect 66626 15750 66638 15802
rect 66690 15750 66702 15802
rect 66754 15750 66766 15802
rect 66818 15750 66830 15802
rect 66882 15750 77924 15802
rect 2024 15728 77924 15750
rect 2024 15258 77924 15280
rect 2024 15206 5794 15258
rect 5846 15206 5858 15258
rect 5910 15206 5922 15258
rect 5974 15206 5986 15258
rect 6038 15206 6050 15258
rect 6102 15206 36514 15258
rect 36566 15206 36578 15258
rect 36630 15206 36642 15258
rect 36694 15206 36706 15258
rect 36758 15206 36770 15258
rect 36822 15206 67234 15258
rect 67286 15206 67298 15258
rect 67350 15206 67362 15258
rect 67414 15206 67426 15258
rect 67478 15206 67490 15258
rect 67542 15206 77924 15258
rect 2024 15184 77924 15206
rect 2024 14714 77924 14736
rect 2024 14662 5134 14714
rect 5186 14662 5198 14714
rect 5250 14662 5262 14714
rect 5314 14662 5326 14714
rect 5378 14662 5390 14714
rect 5442 14662 35854 14714
rect 35906 14662 35918 14714
rect 35970 14662 35982 14714
rect 36034 14662 36046 14714
rect 36098 14662 36110 14714
rect 36162 14662 66574 14714
rect 66626 14662 66638 14714
rect 66690 14662 66702 14714
rect 66754 14662 66766 14714
rect 66818 14662 66830 14714
rect 66882 14662 77924 14714
rect 2024 14640 77924 14662
rect 2024 14170 77924 14192
rect 2024 14118 5794 14170
rect 5846 14118 5858 14170
rect 5910 14118 5922 14170
rect 5974 14118 5986 14170
rect 6038 14118 6050 14170
rect 6102 14118 36514 14170
rect 36566 14118 36578 14170
rect 36630 14118 36642 14170
rect 36694 14118 36706 14170
rect 36758 14118 36770 14170
rect 36822 14118 67234 14170
rect 67286 14118 67298 14170
rect 67350 14118 67362 14170
rect 67414 14118 67426 14170
rect 67478 14118 67490 14170
rect 67542 14118 77924 14170
rect 2024 14096 77924 14118
rect 2024 13626 77924 13648
rect 2024 13574 5134 13626
rect 5186 13574 5198 13626
rect 5250 13574 5262 13626
rect 5314 13574 5326 13626
rect 5378 13574 5390 13626
rect 5442 13574 35854 13626
rect 35906 13574 35918 13626
rect 35970 13574 35982 13626
rect 36034 13574 36046 13626
rect 36098 13574 36110 13626
rect 36162 13574 66574 13626
rect 66626 13574 66638 13626
rect 66690 13574 66702 13626
rect 66754 13574 66766 13626
rect 66818 13574 66830 13626
rect 66882 13574 77924 13626
rect 2024 13552 77924 13574
rect 2024 13082 77924 13104
rect 2024 13030 5794 13082
rect 5846 13030 5858 13082
rect 5910 13030 5922 13082
rect 5974 13030 5986 13082
rect 6038 13030 6050 13082
rect 6102 13030 36514 13082
rect 36566 13030 36578 13082
rect 36630 13030 36642 13082
rect 36694 13030 36706 13082
rect 36758 13030 36770 13082
rect 36822 13030 67234 13082
rect 67286 13030 67298 13082
rect 67350 13030 67362 13082
rect 67414 13030 67426 13082
rect 67478 13030 67490 13082
rect 67542 13030 77924 13082
rect 2024 13008 77924 13030
rect 2024 12538 77924 12560
rect 2024 12486 5134 12538
rect 5186 12486 5198 12538
rect 5250 12486 5262 12538
rect 5314 12486 5326 12538
rect 5378 12486 5390 12538
rect 5442 12486 35854 12538
rect 35906 12486 35918 12538
rect 35970 12486 35982 12538
rect 36034 12486 36046 12538
rect 36098 12486 36110 12538
rect 36162 12486 66574 12538
rect 66626 12486 66638 12538
rect 66690 12486 66702 12538
rect 66754 12486 66766 12538
rect 66818 12486 66830 12538
rect 66882 12486 77924 12538
rect 2024 12464 77924 12486
rect 2024 11994 77924 12016
rect 2024 11942 5794 11994
rect 5846 11942 5858 11994
rect 5910 11942 5922 11994
rect 5974 11942 5986 11994
rect 6038 11942 6050 11994
rect 6102 11942 36514 11994
rect 36566 11942 36578 11994
rect 36630 11942 36642 11994
rect 36694 11942 36706 11994
rect 36758 11942 36770 11994
rect 36822 11942 67234 11994
rect 67286 11942 67298 11994
rect 67350 11942 67362 11994
rect 67414 11942 67426 11994
rect 67478 11942 67490 11994
rect 67542 11942 77924 11994
rect 2024 11920 77924 11942
rect 2024 11450 77924 11472
rect 2024 11398 5134 11450
rect 5186 11398 5198 11450
rect 5250 11398 5262 11450
rect 5314 11398 5326 11450
rect 5378 11398 5390 11450
rect 5442 11398 35854 11450
rect 35906 11398 35918 11450
rect 35970 11398 35982 11450
rect 36034 11398 36046 11450
rect 36098 11398 36110 11450
rect 36162 11398 66574 11450
rect 66626 11398 66638 11450
rect 66690 11398 66702 11450
rect 66754 11398 66766 11450
rect 66818 11398 66830 11450
rect 66882 11398 77924 11450
rect 2024 11376 77924 11398
rect 2024 10906 77924 10928
rect 2024 10854 5794 10906
rect 5846 10854 5858 10906
rect 5910 10854 5922 10906
rect 5974 10854 5986 10906
rect 6038 10854 6050 10906
rect 6102 10854 36514 10906
rect 36566 10854 36578 10906
rect 36630 10854 36642 10906
rect 36694 10854 36706 10906
rect 36758 10854 36770 10906
rect 36822 10854 67234 10906
rect 67286 10854 67298 10906
rect 67350 10854 67362 10906
rect 67414 10854 67426 10906
rect 67478 10854 67490 10906
rect 67542 10854 77924 10906
rect 2024 10832 77924 10854
rect 2024 10362 77924 10384
rect 2024 10310 5134 10362
rect 5186 10310 5198 10362
rect 5250 10310 5262 10362
rect 5314 10310 5326 10362
rect 5378 10310 5390 10362
rect 5442 10310 35854 10362
rect 35906 10310 35918 10362
rect 35970 10310 35982 10362
rect 36034 10310 36046 10362
rect 36098 10310 36110 10362
rect 36162 10310 66574 10362
rect 66626 10310 66638 10362
rect 66690 10310 66702 10362
rect 66754 10310 66766 10362
rect 66818 10310 66830 10362
rect 66882 10310 77924 10362
rect 2024 10288 77924 10310
rect 2024 9818 77924 9840
rect 2024 9766 5794 9818
rect 5846 9766 5858 9818
rect 5910 9766 5922 9818
rect 5974 9766 5986 9818
rect 6038 9766 6050 9818
rect 6102 9766 36514 9818
rect 36566 9766 36578 9818
rect 36630 9766 36642 9818
rect 36694 9766 36706 9818
rect 36758 9766 36770 9818
rect 36822 9766 67234 9818
rect 67286 9766 67298 9818
rect 67350 9766 67362 9818
rect 67414 9766 67426 9818
rect 67478 9766 67490 9818
rect 67542 9766 77924 9818
rect 2024 9744 77924 9766
rect 2024 9274 77924 9296
rect 2024 9222 5134 9274
rect 5186 9222 5198 9274
rect 5250 9222 5262 9274
rect 5314 9222 5326 9274
rect 5378 9222 5390 9274
rect 5442 9222 35854 9274
rect 35906 9222 35918 9274
rect 35970 9222 35982 9274
rect 36034 9222 36046 9274
rect 36098 9222 36110 9274
rect 36162 9222 66574 9274
rect 66626 9222 66638 9274
rect 66690 9222 66702 9274
rect 66754 9222 66766 9274
rect 66818 9222 66830 9274
rect 66882 9222 77924 9274
rect 2024 9200 77924 9222
rect 2024 8730 77924 8752
rect 2024 8678 5794 8730
rect 5846 8678 5858 8730
rect 5910 8678 5922 8730
rect 5974 8678 5986 8730
rect 6038 8678 6050 8730
rect 6102 8678 36514 8730
rect 36566 8678 36578 8730
rect 36630 8678 36642 8730
rect 36694 8678 36706 8730
rect 36758 8678 36770 8730
rect 36822 8678 67234 8730
rect 67286 8678 67298 8730
rect 67350 8678 67362 8730
rect 67414 8678 67426 8730
rect 67478 8678 67490 8730
rect 67542 8678 77924 8730
rect 2024 8656 77924 8678
rect 2024 8186 77924 8208
rect 2024 8134 5134 8186
rect 5186 8134 5198 8186
rect 5250 8134 5262 8186
rect 5314 8134 5326 8186
rect 5378 8134 5390 8186
rect 5442 8134 35854 8186
rect 35906 8134 35918 8186
rect 35970 8134 35982 8186
rect 36034 8134 36046 8186
rect 36098 8134 36110 8186
rect 36162 8134 66574 8186
rect 66626 8134 66638 8186
rect 66690 8134 66702 8186
rect 66754 8134 66766 8186
rect 66818 8134 66830 8186
rect 66882 8134 77924 8186
rect 2024 8112 77924 8134
rect 2024 7642 77924 7664
rect 2024 7590 5794 7642
rect 5846 7590 5858 7642
rect 5910 7590 5922 7642
rect 5974 7590 5986 7642
rect 6038 7590 6050 7642
rect 6102 7590 36514 7642
rect 36566 7590 36578 7642
rect 36630 7590 36642 7642
rect 36694 7590 36706 7642
rect 36758 7590 36770 7642
rect 36822 7590 67234 7642
rect 67286 7590 67298 7642
rect 67350 7590 67362 7642
rect 67414 7590 67426 7642
rect 67478 7590 67490 7642
rect 67542 7590 77924 7642
rect 2024 7568 77924 7590
rect 2024 7098 77924 7120
rect 2024 7046 5134 7098
rect 5186 7046 5198 7098
rect 5250 7046 5262 7098
rect 5314 7046 5326 7098
rect 5378 7046 5390 7098
rect 5442 7046 35854 7098
rect 35906 7046 35918 7098
rect 35970 7046 35982 7098
rect 36034 7046 36046 7098
rect 36098 7046 36110 7098
rect 36162 7046 66574 7098
rect 66626 7046 66638 7098
rect 66690 7046 66702 7098
rect 66754 7046 66766 7098
rect 66818 7046 66830 7098
rect 66882 7046 77924 7098
rect 2024 7024 77924 7046
rect 2024 6554 77924 6576
rect 2024 6502 5794 6554
rect 5846 6502 5858 6554
rect 5910 6502 5922 6554
rect 5974 6502 5986 6554
rect 6038 6502 6050 6554
rect 6102 6502 36514 6554
rect 36566 6502 36578 6554
rect 36630 6502 36642 6554
rect 36694 6502 36706 6554
rect 36758 6502 36770 6554
rect 36822 6502 67234 6554
rect 67286 6502 67298 6554
rect 67350 6502 67362 6554
rect 67414 6502 67426 6554
rect 67478 6502 67490 6554
rect 67542 6502 77924 6554
rect 2024 6480 77924 6502
rect 2024 6010 77924 6032
rect 2024 5958 5134 6010
rect 5186 5958 5198 6010
rect 5250 5958 5262 6010
rect 5314 5958 5326 6010
rect 5378 5958 5390 6010
rect 5442 5958 35854 6010
rect 35906 5958 35918 6010
rect 35970 5958 35982 6010
rect 36034 5958 36046 6010
rect 36098 5958 36110 6010
rect 36162 5958 66574 6010
rect 66626 5958 66638 6010
rect 66690 5958 66702 6010
rect 66754 5958 66766 6010
rect 66818 5958 66830 6010
rect 66882 5958 77924 6010
rect 2024 5936 77924 5958
rect 2024 5466 77924 5488
rect 2024 5414 5794 5466
rect 5846 5414 5858 5466
rect 5910 5414 5922 5466
rect 5974 5414 5986 5466
rect 6038 5414 6050 5466
rect 6102 5414 36514 5466
rect 36566 5414 36578 5466
rect 36630 5414 36642 5466
rect 36694 5414 36706 5466
rect 36758 5414 36770 5466
rect 36822 5414 67234 5466
rect 67286 5414 67298 5466
rect 67350 5414 67362 5466
rect 67414 5414 67426 5466
rect 67478 5414 67490 5466
rect 67542 5414 77924 5466
rect 2024 5392 77924 5414
rect 2024 4922 77924 4944
rect 2024 4870 5134 4922
rect 5186 4870 5198 4922
rect 5250 4870 5262 4922
rect 5314 4870 5326 4922
rect 5378 4870 5390 4922
rect 5442 4870 35854 4922
rect 35906 4870 35918 4922
rect 35970 4870 35982 4922
rect 36034 4870 36046 4922
rect 36098 4870 36110 4922
rect 36162 4870 66574 4922
rect 66626 4870 66638 4922
rect 66690 4870 66702 4922
rect 66754 4870 66766 4922
rect 66818 4870 66830 4922
rect 66882 4870 77924 4922
rect 2024 4848 77924 4870
rect 2024 4378 77924 4400
rect 2024 4326 5794 4378
rect 5846 4326 5858 4378
rect 5910 4326 5922 4378
rect 5974 4326 5986 4378
rect 6038 4326 6050 4378
rect 6102 4326 36514 4378
rect 36566 4326 36578 4378
rect 36630 4326 36642 4378
rect 36694 4326 36706 4378
rect 36758 4326 36770 4378
rect 36822 4326 67234 4378
rect 67286 4326 67298 4378
rect 67350 4326 67362 4378
rect 67414 4326 67426 4378
rect 67478 4326 67490 4378
rect 67542 4326 77924 4378
rect 2024 4304 77924 4326
rect 2024 3834 77924 3856
rect 2024 3782 5134 3834
rect 5186 3782 5198 3834
rect 5250 3782 5262 3834
rect 5314 3782 5326 3834
rect 5378 3782 5390 3834
rect 5442 3782 35854 3834
rect 35906 3782 35918 3834
rect 35970 3782 35982 3834
rect 36034 3782 36046 3834
rect 36098 3782 36110 3834
rect 36162 3782 66574 3834
rect 66626 3782 66638 3834
rect 66690 3782 66702 3834
rect 66754 3782 66766 3834
rect 66818 3782 66830 3834
rect 66882 3782 77924 3834
rect 2024 3760 77924 3782
rect 2024 3290 77924 3312
rect 2024 3238 5794 3290
rect 5846 3238 5858 3290
rect 5910 3238 5922 3290
rect 5974 3238 5986 3290
rect 6038 3238 6050 3290
rect 6102 3238 36514 3290
rect 36566 3238 36578 3290
rect 36630 3238 36642 3290
rect 36694 3238 36706 3290
rect 36758 3238 36770 3290
rect 36822 3238 67234 3290
rect 67286 3238 67298 3290
rect 67350 3238 67362 3290
rect 67414 3238 67426 3290
rect 67478 3238 67490 3290
rect 67542 3238 77924 3290
rect 2024 3216 77924 3238
rect 2024 2746 77924 2768
rect 2024 2694 5134 2746
rect 5186 2694 5198 2746
rect 5250 2694 5262 2746
rect 5314 2694 5326 2746
rect 5378 2694 5390 2746
rect 5442 2694 35854 2746
rect 35906 2694 35918 2746
rect 35970 2694 35982 2746
rect 36034 2694 36046 2746
rect 36098 2694 36110 2746
rect 36162 2694 66574 2746
rect 66626 2694 66638 2746
rect 66690 2694 66702 2746
rect 66754 2694 66766 2746
rect 66818 2694 66830 2746
rect 66882 2694 77924 2746
rect 2024 2672 77924 2694
rect 22554 2388 22560 2440
rect 22612 2428 22618 2440
rect 22741 2431 22799 2437
rect 22741 2428 22753 2431
rect 22612 2400 22753 2428
rect 22612 2388 22618 2400
rect 22741 2397 22753 2400
rect 22787 2397 22799 2431
rect 22741 2391 22799 2397
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23293 2431 23351 2437
rect 23293 2428 23305 2431
rect 23256 2400 23305 2428
rect 23256 2388 23262 2400
rect 23293 2397 23305 2400
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33560 2400 33609 2428
rect 33560 2388 33566 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 33597 2391 33655 2397
rect 41874 2388 41880 2440
rect 41932 2428 41938 2440
rect 41969 2431 42027 2437
rect 41969 2428 41981 2431
rect 41932 2400 41981 2428
rect 41932 2388 41938 2400
rect 41969 2397 41981 2400
rect 42015 2397 42027 2431
rect 41969 2391 42027 2397
rect 42518 2388 42524 2440
rect 42576 2428 42582 2440
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 42576 2400 42625 2428
rect 42576 2388 42582 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 42613 2391 42671 2397
rect 44450 2388 44456 2440
rect 44508 2428 44514 2440
rect 44545 2431 44603 2437
rect 44545 2428 44557 2431
rect 44508 2400 44557 2428
rect 44508 2388 44514 2400
rect 44545 2397 44557 2400
rect 44591 2397 44603 2431
rect 44545 2391 44603 2397
rect 52178 2388 52184 2440
rect 52236 2428 52242 2440
rect 52273 2431 52331 2437
rect 52273 2428 52285 2431
rect 52236 2400 52285 2428
rect 52236 2388 52242 2400
rect 52273 2397 52285 2400
rect 52319 2397 52331 2431
rect 52273 2391 52331 2397
rect 57974 2388 57980 2440
rect 58032 2428 58038 2440
rect 58069 2431 58127 2437
rect 58069 2428 58081 2431
rect 58032 2400 58081 2428
rect 58032 2388 58038 2400
rect 58069 2397 58081 2400
rect 58115 2397 58127 2431
rect 58069 2391 58127 2397
rect 59262 2388 59268 2440
rect 59320 2428 59326 2440
rect 59357 2431 59415 2437
rect 59357 2428 59369 2431
rect 59320 2400 59369 2428
rect 59320 2388 59326 2400
rect 59357 2397 59369 2400
rect 59403 2397 59415 2431
rect 59357 2391 59415 2397
rect 2024 2202 77924 2224
rect 2024 2150 5794 2202
rect 5846 2150 5858 2202
rect 5910 2150 5922 2202
rect 5974 2150 5986 2202
rect 6038 2150 6050 2202
rect 6102 2150 36514 2202
rect 36566 2150 36578 2202
rect 36630 2150 36642 2202
rect 36694 2150 36706 2202
rect 36758 2150 36770 2202
rect 36822 2150 67234 2202
rect 67286 2150 67298 2202
rect 67350 2150 67362 2202
rect 67414 2150 67426 2202
rect 67478 2150 67490 2202
rect 67542 2150 77924 2202
rect 2024 2128 77924 2150
<< via1 >>
rect 5134 77766 5186 77818
rect 5198 77766 5250 77818
rect 5262 77766 5314 77818
rect 5326 77766 5378 77818
rect 5390 77766 5442 77818
rect 35854 77766 35906 77818
rect 35918 77766 35970 77818
rect 35982 77766 36034 77818
rect 36046 77766 36098 77818
rect 36110 77766 36162 77818
rect 66574 77766 66626 77818
rect 66638 77766 66690 77818
rect 66702 77766 66754 77818
rect 66766 77766 66818 77818
rect 66830 77766 66882 77818
rect 23848 77664 23900 77716
rect 32864 77664 32916 77716
rect 39948 77664 40000 77716
rect 41880 77664 41932 77716
rect 49608 77664 49660 77716
rect 54116 77664 54168 77716
rect 58624 77664 58676 77716
rect 5794 77222 5846 77274
rect 5858 77222 5910 77274
rect 5922 77222 5974 77274
rect 5986 77222 6038 77274
rect 6050 77222 6102 77274
rect 36514 77222 36566 77274
rect 36578 77222 36630 77274
rect 36642 77222 36694 77274
rect 36706 77222 36758 77274
rect 36770 77222 36822 77274
rect 67234 77222 67286 77274
rect 67298 77222 67350 77274
rect 67362 77222 67414 77274
rect 67426 77222 67478 77274
rect 67490 77222 67542 77274
rect 5134 76678 5186 76730
rect 5198 76678 5250 76730
rect 5262 76678 5314 76730
rect 5326 76678 5378 76730
rect 5390 76678 5442 76730
rect 35854 76678 35906 76730
rect 35918 76678 35970 76730
rect 35982 76678 36034 76730
rect 36046 76678 36098 76730
rect 36110 76678 36162 76730
rect 66574 76678 66626 76730
rect 66638 76678 66690 76730
rect 66702 76678 66754 76730
rect 66766 76678 66818 76730
rect 66830 76678 66882 76730
rect 5794 76134 5846 76186
rect 5858 76134 5910 76186
rect 5922 76134 5974 76186
rect 5986 76134 6038 76186
rect 6050 76134 6102 76186
rect 36514 76134 36566 76186
rect 36578 76134 36630 76186
rect 36642 76134 36694 76186
rect 36706 76134 36758 76186
rect 36770 76134 36822 76186
rect 67234 76134 67286 76186
rect 67298 76134 67350 76186
rect 67362 76134 67414 76186
rect 67426 76134 67478 76186
rect 67490 76134 67542 76186
rect 5134 75590 5186 75642
rect 5198 75590 5250 75642
rect 5262 75590 5314 75642
rect 5326 75590 5378 75642
rect 5390 75590 5442 75642
rect 35854 75590 35906 75642
rect 35918 75590 35970 75642
rect 35982 75590 36034 75642
rect 36046 75590 36098 75642
rect 36110 75590 36162 75642
rect 66574 75590 66626 75642
rect 66638 75590 66690 75642
rect 66702 75590 66754 75642
rect 66766 75590 66818 75642
rect 66830 75590 66882 75642
rect 5794 75046 5846 75098
rect 5858 75046 5910 75098
rect 5922 75046 5974 75098
rect 5986 75046 6038 75098
rect 6050 75046 6102 75098
rect 36514 75046 36566 75098
rect 36578 75046 36630 75098
rect 36642 75046 36694 75098
rect 36706 75046 36758 75098
rect 36770 75046 36822 75098
rect 67234 75046 67286 75098
rect 67298 75046 67350 75098
rect 67362 75046 67414 75098
rect 67426 75046 67478 75098
rect 67490 75046 67542 75098
rect 5134 74502 5186 74554
rect 5198 74502 5250 74554
rect 5262 74502 5314 74554
rect 5326 74502 5378 74554
rect 5390 74502 5442 74554
rect 35854 74502 35906 74554
rect 35918 74502 35970 74554
rect 35982 74502 36034 74554
rect 36046 74502 36098 74554
rect 36110 74502 36162 74554
rect 66574 74502 66626 74554
rect 66638 74502 66690 74554
rect 66702 74502 66754 74554
rect 66766 74502 66818 74554
rect 66830 74502 66882 74554
rect 5794 73958 5846 74010
rect 5858 73958 5910 74010
rect 5922 73958 5974 74010
rect 5986 73958 6038 74010
rect 6050 73958 6102 74010
rect 36514 73958 36566 74010
rect 36578 73958 36630 74010
rect 36642 73958 36694 74010
rect 36706 73958 36758 74010
rect 36770 73958 36822 74010
rect 67234 73958 67286 74010
rect 67298 73958 67350 74010
rect 67362 73958 67414 74010
rect 67426 73958 67478 74010
rect 67490 73958 67542 74010
rect 5134 73414 5186 73466
rect 5198 73414 5250 73466
rect 5262 73414 5314 73466
rect 5326 73414 5378 73466
rect 5390 73414 5442 73466
rect 35854 73414 35906 73466
rect 35918 73414 35970 73466
rect 35982 73414 36034 73466
rect 36046 73414 36098 73466
rect 36110 73414 36162 73466
rect 66574 73414 66626 73466
rect 66638 73414 66690 73466
rect 66702 73414 66754 73466
rect 66766 73414 66818 73466
rect 66830 73414 66882 73466
rect 5794 72870 5846 72922
rect 5858 72870 5910 72922
rect 5922 72870 5974 72922
rect 5986 72870 6038 72922
rect 6050 72870 6102 72922
rect 36514 72870 36566 72922
rect 36578 72870 36630 72922
rect 36642 72870 36694 72922
rect 36706 72870 36758 72922
rect 36770 72870 36822 72922
rect 67234 72870 67286 72922
rect 67298 72870 67350 72922
rect 67362 72870 67414 72922
rect 67426 72870 67478 72922
rect 67490 72870 67542 72922
rect 5134 72326 5186 72378
rect 5198 72326 5250 72378
rect 5262 72326 5314 72378
rect 5326 72326 5378 72378
rect 5390 72326 5442 72378
rect 35854 72326 35906 72378
rect 35918 72326 35970 72378
rect 35982 72326 36034 72378
rect 36046 72326 36098 72378
rect 36110 72326 36162 72378
rect 66574 72326 66626 72378
rect 66638 72326 66690 72378
rect 66702 72326 66754 72378
rect 66766 72326 66818 72378
rect 66830 72326 66882 72378
rect 5794 71782 5846 71834
rect 5858 71782 5910 71834
rect 5922 71782 5974 71834
rect 5986 71782 6038 71834
rect 6050 71782 6102 71834
rect 36514 71782 36566 71834
rect 36578 71782 36630 71834
rect 36642 71782 36694 71834
rect 36706 71782 36758 71834
rect 36770 71782 36822 71834
rect 67234 71782 67286 71834
rect 67298 71782 67350 71834
rect 67362 71782 67414 71834
rect 67426 71782 67478 71834
rect 67490 71782 67542 71834
rect 5134 71238 5186 71290
rect 5198 71238 5250 71290
rect 5262 71238 5314 71290
rect 5326 71238 5378 71290
rect 5390 71238 5442 71290
rect 35854 71238 35906 71290
rect 35918 71238 35970 71290
rect 35982 71238 36034 71290
rect 36046 71238 36098 71290
rect 36110 71238 36162 71290
rect 66574 71238 66626 71290
rect 66638 71238 66690 71290
rect 66702 71238 66754 71290
rect 66766 71238 66818 71290
rect 66830 71238 66882 71290
rect 5794 70694 5846 70746
rect 5858 70694 5910 70746
rect 5922 70694 5974 70746
rect 5986 70694 6038 70746
rect 6050 70694 6102 70746
rect 36514 70694 36566 70746
rect 36578 70694 36630 70746
rect 36642 70694 36694 70746
rect 36706 70694 36758 70746
rect 36770 70694 36822 70746
rect 67234 70694 67286 70746
rect 67298 70694 67350 70746
rect 67362 70694 67414 70746
rect 67426 70694 67478 70746
rect 67490 70694 67542 70746
rect 5134 70150 5186 70202
rect 5198 70150 5250 70202
rect 5262 70150 5314 70202
rect 5326 70150 5378 70202
rect 5390 70150 5442 70202
rect 35854 70150 35906 70202
rect 35918 70150 35970 70202
rect 35982 70150 36034 70202
rect 36046 70150 36098 70202
rect 36110 70150 36162 70202
rect 66574 70150 66626 70202
rect 66638 70150 66690 70202
rect 66702 70150 66754 70202
rect 66766 70150 66818 70202
rect 66830 70150 66882 70202
rect 5794 69606 5846 69658
rect 5858 69606 5910 69658
rect 5922 69606 5974 69658
rect 5986 69606 6038 69658
rect 6050 69606 6102 69658
rect 36514 69606 36566 69658
rect 36578 69606 36630 69658
rect 36642 69606 36694 69658
rect 36706 69606 36758 69658
rect 36770 69606 36822 69658
rect 67234 69606 67286 69658
rect 67298 69606 67350 69658
rect 67362 69606 67414 69658
rect 67426 69606 67478 69658
rect 67490 69606 67542 69658
rect 5134 69062 5186 69114
rect 5198 69062 5250 69114
rect 5262 69062 5314 69114
rect 5326 69062 5378 69114
rect 5390 69062 5442 69114
rect 35854 69062 35906 69114
rect 35918 69062 35970 69114
rect 35982 69062 36034 69114
rect 36046 69062 36098 69114
rect 36110 69062 36162 69114
rect 66574 69062 66626 69114
rect 66638 69062 66690 69114
rect 66702 69062 66754 69114
rect 66766 69062 66818 69114
rect 66830 69062 66882 69114
rect 5794 68518 5846 68570
rect 5858 68518 5910 68570
rect 5922 68518 5974 68570
rect 5986 68518 6038 68570
rect 6050 68518 6102 68570
rect 36514 68518 36566 68570
rect 36578 68518 36630 68570
rect 36642 68518 36694 68570
rect 36706 68518 36758 68570
rect 36770 68518 36822 68570
rect 67234 68518 67286 68570
rect 67298 68518 67350 68570
rect 67362 68518 67414 68570
rect 67426 68518 67478 68570
rect 67490 68518 67542 68570
rect 5134 67974 5186 68026
rect 5198 67974 5250 68026
rect 5262 67974 5314 68026
rect 5326 67974 5378 68026
rect 5390 67974 5442 68026
rect 35854 67974 35906 68026
rect 35918 67974 35970 68026
rect 35982 67974 36034 68026
rect 36046 67974 36098 68026
rect 36110 67974 36162 68026
rect 66574 67974 66626 68026
rect 66638 67974 66690 68026
rect 66702 67974 66754 68026
rect 66766 67974 66818 68026
rect 66830 67974 66882 68026
rect 5794 67430 5846 67482
rect 5858 67430 5910 67482
rect 5922 67430 5974 67482
rect 5986 67430 6038 67482
rect 6050 67430 6102 67482
rect 36514 67430 36566 67482
rect 36578 67430 36630 67482
rect 36642 67430 36694 67482
rect 36706 67430 36758 67482
rect 36770 67430 36822 67482
rect 67234 67430 67286 67482
rect 67298 67430 67350 67482
rect 67362 67430 67414 67482
rect 67426 67430 67478 67482
rect 67490 67430 67542 67482
rect 5134 66886 5186 66938
rect 5198 66886 5250 66938
rect 5262 66886 5314 66938
rect 5326 66886 5378 66938
rect 5390 66886 5442 66938
rect 35854 66886 35906 66938
rect 35918 66886 35970 66938
rect 35982 66886 36034 66938
rect 36046 66886 36098 66938
rect 36110 66886 36162 66938
rect 66574 66886 66626 66938
rect 66638 66886 66690 66938
rect 66702 66886 66754 66938
rect 66766 66886 66818 66938
rect 66830 66886 66882 66938
rect 5794 66342 5846 66394
rect 5858 66342 5910 66394
rect 5922 66342 5974 66394
rect 5986 66342 6038 66394
rect 6050 66342 6102 66394
rect 36514 66342 36566 66394
rect 36578 66342 36630 66394
rect 36642 66342 36694 66394
rect 36706 66342 36758 66394
rect 36770 66342 36822 66394
rect 67234 66342 67286 66394
rect 67298 66342 67350 66394
rect 67362 66342 67414 66394
rect 67426 66342 67478 66394
rect 67490 66342 67542 66394
rect 5134 65798 5186 65850
rect 5198 65798 5250 65850
rect 5262 65798 5314 65850
rect 5326 65798 5378 65850
rect 5390 65798 5442 65850
rect 35854 65798 35906 65850
rect 35918 65798 35970 65850
rect 35982 65798 36034 65850
rect 36046 65798 36098 65850
rect 36110 65798 36162 65850
rect 66574 65798 66626 65850
rect 66638 65798 66690 65850
rect 66702 65798 66754 65850
rect 66766 65798 66818 65850
rect 66830 65798 66882 65850
rect 5794 65254 5846 65306
rect 5858 65254 5910 65306
rect 5922 65254 5974 65306
rect 5986 65254 6038 65306
rect 6050 65254 6102 65306
rect 36514 65254 36566 65306
rect 36578 65254 36630 65306
rect 36642 65254 36694 65306
rect 36706 65254 36758 65306
rect 36770 65254 36822 65306
rect 67234 65254 67286 65306
rect 67298 65254 67350 65306
rect 67362 65254 67414 65306
rect 67426 65254 67478 65306
rect 67490 65254 67542 65306
rect 5134 64710 5186 64762
rect 5198 64710 5250 64762
rect 5262 64710 5314 64762
rect 5326 64710 5378 64762
rect 5390 64710 5442 64762
rect 35854 64710 35906 64762
rect 35918 64710 35970 64762
rect 35982 64710 36034 64762
rect 36046 64710 36098 64762
rect 36110 64710 36162 64762
rect 66574 64710 66626 64762
rect 66638 64710 66690 64762
rect 66702 64710 66754 64762
rect 66766 64710 66818 64762
rect 66830 64710 66882 64762
rect 5794 64166 5846 64218
rect 5858 64166 5910 64218
rect 5922 64166 5974 64218
rect 5986 64166 6038 64218
rect 6050 64166 6102 64218
rect 36514 64166 36566 64218
rect 36578 64166 36630 64218
rect 36642 64166 36694 64218
rect 36706 64166 36758 64218
rect 36770 64166 36822 64218
rect 67234 64166 67286 64218
rect 67298 64166 67350 64218
rect 67362 64166 67414 64218
rect 67426 64166 67478 64218
rect 67490 64166 67542 64218
rect 5134 63622 5186 63674
rect 5198 63622 5250 63674
rect 5262 63622 5314 63674
rect 5326 63622 5378 63674
rect 5390 63622 5442 63674
rect 35854 63622 35906 63674
rect 35918 63622 35970 63674
rect 35982 63622 36034 63674
rect 36046 63622 36098 63674
rect 36110 63622 36162 63674
rect 66574 63622 66626 63674
rect 66638 63622 66690 63674
rect 66702 63622 66754 63674
rect 66766 63622 66818 63674
rect 66830 63622 66882 63674
rect 5794 63078 5846 63130
rect 5858 63078 5910 63130
rect 5922 63078 5974 63130
rect 5986 63078 6038 63130
rect 6050 63078 6102 63130
rect 36514 63078 36566 63130
rect 36578 63078 36630 63130
rect 36642 63078 36694 63130
rect 36706 63078 36758 63130
rect 36770 63078 36822 63130
rect 67234 63078 67286 63130
rect 67298 63078 67350 63130
rect 67362 63078 67414 63130
rect 67426 63078 67478 63130
rect 67490 63078 67542 63130
rect 5134 62534 5186 62586
rect 5198 62534 5250 62586
rect 5262 62534 5314 62586
rect 5326 62534 5378 62586
rect 5390 62534 5442 62586
rect 35854 62534 35906 62586
rect 35918 62534 35970 62586
rect 35982 62534 36034 62586
rect 36046 62534 36098 62586
rect 36110 62534 36162 62586
rect 66574 62534 66626 62586
rect 66638 62534 66690 62586
rect 66702 62534 66754 62586
rect 66766 62534 66818 62586
rect 66830 62534 66882 62586
rect 5794 61990 5846 62042
rect 5858 61990 5910 62042
rect 5922 61990 5974 62042
rect 5986 61990 6038 62042
rect 6050 61990 6102 62042
rect 36514 61990 36566 62042
rect 36578 61990 36630 62042
rect 36642 61990 36694 62042
rect 36706 61990 36758 62042
rect 36770 61990 36822 62042
rect 67234 61990 67286 62042
rect 67298 61990 67350 62042
rect 67362 61990 67414 62042
rect 67426 61990 67478 62042
rect 67490 61990 67542 62042
rect 5134 61446 5186 61498
rect 5198 61446 5250 61498
rect 5262 61446 5314 61498
rect 5326 61446 5378 61498
rect 5390 61446 5442 61498
rect 35854 61446 35906 61498
rect 35918 61446 35970 61498
rect 35982 61446 36034 61498
rect 36046 61446 36098 61498
rect 36110 61446 36162 61498
rect 66574 61446 66626 61498
rect 66638 61446 66690 61498
rect 66702 61446 66754 61498
rect 66766 61446 66818 61498
rect 66830 61446 66882 61498
rect 5794 60902 5846 60954
rect 5858 60902 5910 60954
rect 5922 60902 5974 60954
rect 5986 60902 6038 60954
rect 6050 60902 6102 60954
rect 36514 60902 36566 60954
rect 36578 60902 36630 60954
rect 36642 60902 36694 60954
rect 36706 60902 36758 60954
rect 36770 60902 36822 60954
rect 67234 60902 67286 60954
rect 67298 60902 67350 60954
rect 67362 60902 67414 60954
rect 67426 60902 67478 60954
rect 67490 60902 67542 60954
rect 5134 60358 5186 60410
rect 5198 60358 5250 60410
rect 5262 60358 5314 60410
rect 5326 60358 5378 60410
rect 5390 60358 5442 60410
rect 35854 60358 35906 60410
rect 35918 60358 35970 60410
rect 35982 60358 36034 60410
rect 36046 60358 36098 60410
rect 36110 60358 36162 60410
rect 66574 60358 66626 60410
rect 66638 60358 66690 60410
rect 66702 60358 66754 60410
rect 66766 60358 66818 60410
rect 66830 60358 66882 60410
rect 5794 59814 5846 59866
rect 5858 59814 5910 59866
rect 5922 59814 5974 59866
rect 5986 59814 6038 59866
rect 6050 59814 6102 59866
rect 36514 59814 36566 59866
rect 36578 59814 36630 59866
rect 36642 59814 36694 59866
rect 36706 59814 36758 59866
rect 36770 59814 36822 59866
rect 67234 59814 67286 59866
rect 67298 59814 67350 59866
rect 67362 59814 67414 59866
rect 67426 59814 67478 59866
rect 67490 59814 67542 59866
rect 5134 59270 5186 59322
rect 5198 59270 5250 59322
rect 5262 59270 5314 59322
rect 5326 59270 5378 59322
rect 5390 59270 5442 59322
rect 35854 59270 35906 59322
rect 35918 59270 35970 59322
rect 35982 59270 36034 59322
rect 36046 59270 36098 59322
rect 36110 59270 36162 59322
rect 66574 59270 66626 59322
rect 66638 59270 66690 59322
rect 66702 59270 66754 59322
rect 66766 59270 66818 59322
rect 66830 59270 66882 59322
rect 5794 58726 5846 58778
rect 5858 58726 5910 58778
rect 5922 58726 5974 58778
rect 5986 58726 6038 58778
rect 6050 58726 6102 58778
rect 36514 58726 36566 58778
rect 36578 58726 36630 58778
rect 36642 58726 36694 58778
rect 36706 58726 36758 58778
rect 36770 58726 36822 58778
rect 67234 58726 67286 58778
rect 67298 58726 67350 58778
rect 67362 58726 67414 58778
rect 67426 58726 67478 58778
rect 67490 58726 67542 58778
rect 5134 58182 5186 58234
rect 5198 58182 5250 58234
rect 5262 58182 5314 58234
rect 5326 58182 5378 58234
rect 5390 58182 5442 58234
rect 35854 58182 35906 58234
rect 35918 58182 35970 58234
rect 35982 58182 36034 58234
rect 36046 58182 36098 58234
rect 36110 58182 36162 58234
rect 66574 58182 66626 58234
rect 66638 58182 66690 58234
rect 66702 58182 66754 58234
rect 66766 58182 66818 58234
rect 66830 58182 66882 58234
rect 5794 57638 5846 57690
rect 5858 57638 5910 57690
rect 5922 57638 5974 57690
rect 5986 57638 6038 57690
rect 6050 57638 6102 57690
rect 36514 57638 36566 57690
rect 36578 57638 36630 57690
rect 36642 57638 36694 57690
rect 36706 57638 36758 57690
rect 36770 57638 36822 57690
rect 67234 57638 67286 57690
rect 67298 57638 67350 57690
rect 67362 57638 67414 57690
rect 67426 57638 67478 57690
rect 67490 57638 67542 57690
rect 5134 57094 5186 57146
rect 5198 57094 5250 57146
rect 5262 57094 5314 57146
rect 5326 57094 5378 57146
rect 5390 57094 5442 57146
rect 35854 57094 35906 57146
rect 35918 57094 35970 57146
rect 35982 57094 36034 57146
rect 36046 57094 36098 57146
rect 36110 57094 36162 57146
rect 66574 57094 66626 57146
rect 66638 57094 66690 57146
rect 66702 57094 66754 57146
rect 66766 57094 66818 57146
rect 66830 57094 66882 57146
rect 5794 56550 5846 56602
rect 5858 56550 5910 56602
rect 5922 56550 5974 56602
rect 5986 56550 6038 56602
rect 6050 56550 6102 56602
rect 36514 56550 36566 56602
rect 36578 56550 36630 56602
rect 36642 56550 36694 56602
rect 36706 56550 36758 56602
rect 36770 56550 36822 56602
rect 67234 56550 67286 56602
rect 67298 56550 67350 56602
rect 67362 56550 67414 56602
rect 67426 56550 67478 56602
rect 67490 56550 67542 56602
rect 5134 56006 5186 56058
rect 5198 56006 5250 56058
rect 5262 56006 5314 56058
rect 5326 56006 5378 56058
rect 5390 56006 5442 56058
rect 35854 56006 35906 56058
rect 35918 56006 35970 56058
rect 35982 56006 36034 56058
rect 36046 56006 36098 56058
rect 36110 56006 36162 56058
rect 66574 56006 66626 56058
rect 66638 56006 66690 56058
rect 66702 56006 66754 56058
rect 66766 56006 66818 56058
rect 66830 56006 66882 56058
rect 5794 55462 5846 55514
rect 5858 55462 5910 55514
rect 5922 55462 5974 55514
rect 5986 55462 6038 55514
rect 6050 55462 6102 55514
rect 36514 55462 36566 55514
rect 36578 55462 36630 55514
rect 36642 55462 36694 55514
rect 36706 55462 36758 55514
rect 36770 55462 36822 55514
rect 67234 55462 67286 55514
rect 67298 55462 67350 55514
rect 67362 55462 67414 55514
rect 67426 55462 67478 55514
rect 67490 55462 67542 55514
rect 5134 54918 5186 54970
rect 5198 54918 5250 54970
rect 5262 54918 5314 54970
rect 5326 54918 5378 54970
rect 5390 54918 5442 54970
rect 35854 54918 35906 54970
rect 35918 54918 35970 54970
rect 35982 54918 36034 54970
rect 36046 54918 36098 54970
rect 36110 54918 36162 54970
rect 66574 54918 66626 54970
rect 66638 54918 66690 54970
rect 66702 54918 66754 54970
rect 66766 54918 66818 54970
rect 66830 54918 66882 54970
rect 5794 54374 5846 54426
rect 5858 54374 5910 54426
rect 5922 54374 5974 54426
rect 5986 54374 6038 54426
rect 6050 54374 6102 54426
rect 36514 54374 36566 54426
rect 36578 54374 36630 54426
rect 36642 54374 36694 54426
rect 36706 54374 36758 54426
rect 36770 54374 36822 54426
rect 67234 54374 67286 54426
rect 67298 54374 67350 54426
rect 67362 54374 67414 54426
rect 67426 54374 67478 54426
rect 67490 54374 67542 54426
rect 5134 53830 5186 53882
rect 5198 53830 5250 53882
rect 5262 53830 5314 53882
rect 5326 53830 5378 53882
rect 5390 53830 5442 53882
rect 35854 53830 35906 53882
rect 35918 53830 35970 53882
rect 35982 53830 36034 53882
rect 36046 53830 36098 53882
rect 36110 53830 36162 53882
rect 66574 53830 66626 53882
rect 66638 53830 66690 53882
rect 66702 53830 66754 53882
rect 66766 53830 66818 53882
rect 66830 53830 66882 53882
rect 5794 53286 5846 53338
rect 5858 53286 5910 53338
rect 5922 53286 5974 53338
rect 5986 53286 6038 53338
rect 6050 53286 6102 53338
rect 36514 53286 36566 53338
rect 36578 53286 36630 53338
rect 36642 53286 36694 53338
rect 36706 53286 36758 53338
rect 36770 53286 36822 53338
rect 67234 53286 67286 53338
rect 67298 53286 67350 53338
rect 67362 53286 67414 53338
rect 67426 53286 67478 53338
rect 67490 53286 67542 53338
rect 5134 52742 5186 52794
rect 5198 52742 5250 52794
rect 5262 52742 5314 52794
rect 5326 52742 5378 52794
rect 5390 52742 5442 52794
rect 35854 52742 35906 52794
rect 35918 52742 35970 52794
rect 35982 52742 36034 52794
rect 36046 52742 36098 52794
rect 36110 52742 36162 52794
rect 66574 52742 66626 52794
rect 66638 52742 66690 52794
rect 66702 52742 66754 52794
rect 66766 52742 66818 52794
rect 66830 52742 66882 52794
rect 5794 52198 5846 52250
rect 5858 52198 5910 52250
rect 5922 52198 5974 52250
rect 5986 52198 6038 52250
rect 6050 52198 6102 52250
rect 36514 52198 36566 52250
rect 36578 52198 36630 52250
rect 36642 52198 36694 52250
rect 36706 52198 36758 52250
rect 36770 52198 36822 52250
rect 67234 52198 67286 52250
rect 67298 52198 67350 52250
rect 67362 52198 67414 52250
rect 67426 52198 67478 52250
rect 67490 52198 67542 52250
rect 77576 51799 77628 51808
rect 77576 51765 77585 51799
rect 77585 51765 77619 51799
rect 77619 51765 77628 51799
rect 77576 51756 77628 51765
rect 5134 51654 5186 51706
rect 5198 51654 5250 51706
rect 5262 51654 5314 51706
rect 5326 51654 5378 51706
rect 5390 51654 5442 51706
rect 35854 51654 35906 51706
rect 35918 51654 35970 51706
rect 35982 51654 36034 51706
rect 36046 51654 36098 51706
rect 36110 51654 36162 51706
rect 66574 51654 66626 51706
rect 66638 51654 66690 51706
rect 66702 51654 66754 51706
rect 66766 51654 66818 51706
rect 66830 51654 66882 51706
rect 5794 51110 5846 51162
rect 5858 51110 5910 51162
rect 5922 51110 5974 51162
rect 5986 51110 6038 51162
rect 6050 51110 6102 51162
rect 36514 51110 36566 51162
rect 36578 51110 36630 51162
rect 36642 51110 36694 51162
rect 36706 51110 36758 51162
rect 36770 51110 36822 51162
rect 67234 51110 67286 51162
rect 67298 51110 67350 51162
rect 67362 51110 67414 51162
rect 67426 51110 67478 51162
rect 67490 51110 67542 51162
rect 5134 50566 5186 50618
rect 5198 50566 5250 50618
rect 5262 50566 5314 50618
rect 5326 50566 5378 50618
rect 5390 50566 5442 50618
rect 35854 50566 35906 50618
rect 35918 50566 35970 50618
rect 35982 50566 36034 50618
rect 36046 50566 36098 50618
rect 36110 50566 36162 50618
rect 66574 50566 66626 50618
rect 66638 50566 66690 50618
rect 66702 50566 66754 50618
rect 66766 50566 66818 50618
rect 66830 50566 66882 50618
rect 5794 50022 5846 50074
rect 5858 50022 5910 50074
rect 5922 50022 5974 50074
rect 5986 50022 6038 50074
rect 6050 50022 6102 50074
rect 36514 50022 36566 50074
rect 36578 50022 36630 50074
rect 36642 50022 36694 50074
rect 36706 50022 36758 50074
rect 36770 50022 36822 50074
rect 67234 50022 67286 50074
rect 67298 50022 67350 50074
rect 67362 50022 67414 50074
rect 67426 50022 67478 50074
rect 67490 50022 67542 50074
rect 77576 49759 77628 49768
rect 77576 49725 77585 49759
rect 77585 49725 77619 49759
rect 77619 49725 77628 49759
rect 77576 49716 77628 49725
rect 5134 49478 5186 49530
rect 5198 49478 5250 49530
rect 5262 49478 5314 49530
rect 5326 49478 5378 49530
rect 5390 49478 5442 49530
rect 35854 49478 35906 49530
rect 35918 49478 35970 49530
rect 35982 49478 36034 49530
rect 36046 49478 36098 49530
rect 36110 49478 36162 49530
rect 66574 49478 66626 49530
rect 66638 49478 66690 49530
rect 66702 49478 66754 49530
rect 66766 49478 66818 49530
rect 66830 49478 66882 49530
rect 5794 48934 5846 48986
rect 5858 48934 5910 48986
rect 5922 48934 5974 48986
rect 5986 48934 6038 48986
rect 6050 48934 6102 48986
rect 36514 48934 36566 48986
rect 36578 48934 36630 48986
rect 36642 48934 36694 48986
rect 36706 48934 36758 48986
rect 36770 48934 36822 48986
rect 67234 48934 67286 48986
rect 67298 48934 67350 48986
rect 67362 48934 67414 48986
rect 67426 48934 67478 48986
rect 67490 48934 67542 48986
rect 5134 48390 5186 48442
rect 5198 48390 5250 48442
rect 5262 48390 5314 48442
rect 5326 48390 5378 48442
rect 5390 48390 5442 48442
rect 35854 48390 35906 48442
rect 35918 48390 35970 48442
rect 35982 48390 36034 48442
rect 36046 48390 36098 48442
rect 36110 48390 36162 48442
rect 66574 48390 66626 48442
rect 66638 48390 66690 48442
rect 66702 48390 66754 48442
rect 66766 48390 66818 48442
rect 66830 48390 66882 48442
rect 5794 47846 5846 47898
rect 5858 47846 5910 47898
rect 5922 47846 5974 47898
rect 5986 47846 6038 47898
rect 6050 47846 6102 47898
rect 36514 47846 36566 47898
rect 36578 47846 36630 47898
rect 36642 47846 36694 47898
rect 36706 47846 36758 47898
rect 36770 47846 36822 47898
rect 67234 47846 67286 47898
rect 67298 47846 67350 47898
rect 67362 47846 67414 47898
rect 67426 47846 67478 47898
rect 67490 47846 67542 47898
rect 5134 47302 5186 47354
rect 5198 47302 5250 47354
rect 5262 47302 5314 47354
rect 5326 47302 5378 47354
rect 5390 47302 5442 47354
rect 35854 47302 35906 47354
rect 35918 47302 35970 47354
rect 35982 47302 36034 47354
rect 36046 47302 36098 47354
rect 36110 47302 36162 47354
rect 66574 47302 66626 47354
rect 66638 47302 66690 47354
rect 66702 47302 66754 47354
rect 66766 47302 66818 47354
rect 66830 47302 66882 47354
rect 5794 46758 5846 46810
rect 5858 46758 5910 46810
rect 5922 46758 5974 46810
rect 5986 46758 6038 46810
rect 6050 46758 6102 46810
rect 36514 46758 36566 46810
rect 36578 46758 36630 46810
rect 36642 46758 36694 46810
rect 36706 46758 36758 46810
rect 36770 46758 36822 46810
rect 67234 46758 67286 46810
rect 67298 46758 67350 46810
rect 67362 46758 67414 46810
rect 67426 46758 67478 46810
rect 67490 46758 67542 46810
rect 5134 46214 5186 46266
rect 5198 46214 5250 46266
rect 5262 46214 5314 46266
rect 5326 46214 5378 46266
rect 5390 46214 5442 46266
rect 35854 46214 35906 46266
rect 35918 46214 35970 46266
rect 35982 46214 36034 46266
rect 36046 46214 36098 46266
rect 36110 46214 36162 46266
rect 66574 46214 66626 46266
rect 66638 46214 66690 46266
rect 66702 46214 66754 46266
rect 66766 46214 66818 46266
rect 66830 46214 66882 46266
rect 5794 45670 5846 45722
rect 5858 45670 5910 45722
rect 5922 45670 5974 45722
rect 5986 45670 6038 45722
rect 6050 45670 6102 45722
rect 36514 45670 36566 45722
rect 36578 45670 36630 45722
rect 36642 45670 36694 45722
rect 36706 45670 36758 45722
rect 36770 45670 36822 45722
rect 67234 45670 67286 45722
rect 67298 45670 67350 45722
rect 67362 45670 67414 45722
rect 67426 45670 67478 45722
rect 67490 45670 67542 45722
rect 5134 45126 5186 45178
rect 5198 45126 5250 45178
rect 5262 45126 5314 45178
rect 5326 45126 5378 45178
rect 5390 45126 5442 45178
rect 35854 45126 35906 45178
rect 35918 45126 35970 45178
rect 35982 45126 36034 45178
rect 36046 45126 36098 45178
rect 36110 45126 36162 45178
rect 66574 45126 66626 45178
rect 66638 45126 66690 45178
rect 66702 45126 66754 45178
rect 66766 45126 66818 45178
rect 66830 45126 66882 45178
rect 5794 44582 5846 44634
rect 5858 44582 5910 44634
rect 5922 44582 5974 44634
rect 5986 44582 6038 44634
rect 6050 44582 6102 44634
rect 36514 44582 36566 44634
rect 36578 44582 36630 44634
rect 36642 44582 36694 44634
rect 36706 44582 36758 44634
rect 36770 44582 36822 44634
rect 67234 44582 67286 44634
rect 67298 44582 67350 44634
rect 67362 44582 67414 44634
rect 67426 44582 67478 44634
rect 67490 44582 67542 44634
rect 5134 44038 5186 44090
rect 5198 44038 5250 44090
rect 5262 44038 5314 44090
rect 5326 44038 5378 44090
rect 5390 44038 5442 44090
rect 35854 44038 35906 44090
rect 35918 44038 35970 44090
rect 35982 44038 36034 44090
rect 36046 44038 36098 44090
rect 36110 44038 36162 44090
rect 66574 44038 66626 44090
rect 66638 44038 66690 44090
rect 66702 44038 66754 44090
rect 66766 44038 66818 44090
rect 66830 44038 66882 44090
rect 64880 43843 64932 43852
rect 64880 43809 64889 43843
rect 64889 43809 64923 43843
rect 64923 43809 64932 43843
rect 64880 43800 64932 43809
rect 66904 43732 66956 43784
rect 65432 43596 65484 43648
rect 5794 43494 5846 43546
rect 5858 43494 5910 43546
rect 5922 43494 5974 43546
rect 5986 43494 6038 43546
rect 6050 43494 6102 43546
rect 36514 43494 36566 43546
rect 36578 43494 36630 43546
rect 36642 43494 36694 43546
rect 36706 43494 36758 43546
rect 36770 43494 36822 43546
rect 67234 43494 67286 43546
rect 67298 43494 67350 43546
rect 67362 43494 67414 43546
rect 67426 43494 67478 43546
rect 67490 43494 67542 43546
rect 66260 43392 66312 43444
rect 66904 43435 66956 43444
rect 66904 43401 66913 43435
rect 66913 43401 66947 43435
rect 66947 43401 66956 43435
rect 66904 43392 66956 43401
rect 65432 43367 65484 43376
rect 65432 43333 65441 43367
rect 65441 43333 65475 43367
rect 65475 43333 65484 43367
rect 65432 43324 65484 43333
rect 65156 43231 65208 43240
rect 65156 43197 65165 43231
rect 65165 43197 65199 43231
rect 65199 43197 65208 43231
rect 65156 43188 65208 43197
rect 67088 43188 67140 43240
rect 5134 42950 5186 43002
rect 5198 42950 5250 43002
rect 5262 42950 5314 43002
rect 5326 42950 5378 43002
rect 5390 42950 5442 43002
rect 35854 42950 35906 43002
rect 35918 42950 35970 43002
rect 35982 42950 36034 43002
rect 36046 42950 36098 43002
rect 36110 42950 36162 43002
rect 66574 42950 66626 43002
rect 66638 42950 66690 43002
rect 66702 42950 66754 43002
rect 66766 42950 66818 43002
rect 66830 42950 66882 43002
rect 60004 42712 60056 42764
rect 57612 42687 57664 42696
rect 57612 42653 57621 42687
rect 57621 42653 57655 42687
rect 57655 42653 57664 42687
rect 57612 42644 57664 42653
rect 57980 42576 58032 42628
rect 58900 42576 58952 42628
rect 59544 42551 59596 42560
rect 59544 42517 59553 42551
rect 59553 42517 59587 42551
rect 59587 42517 59596 42551
rect 59544 42508 59596 42517
rect 5794 42406 5846 42458
rect 5858 42406 5910 42458
rect 5922 42406 5974 42458
rect 5986 42406 6038 42458
rect 6050 42406 6102 42458
rect 36514 42406 36566 42458
rect 36578 42406 36630 42458
rect 36642 42406 36694 42458
rect 36706 42406 36758 42458
rect 36770 42406 36822 42458
rect 67234 42406 67286 42458
rect 67298 42406 67350 42458
rect 67362 42406 67414 42458
rect 67426 42406 67478 42458
rect 67490 42406 67542 42458
rect 57980 42304 58032 42356
rect 58900 42347 58952 42356
rect 58900 42313 58909 42347
rect 58909 42313 58943 42347
rect 58943 42313 58952 42347
rect 58900 42304 58952 42313
rect 59544 42236 59596 42288
rect 58992 42211 59044 42220
rect 58992 42177 59001 42211
rect 59001 42177 59035 42211
rect 59035 42177 59044 42211
rect 58992 42168 59044 42177
rect 5134 41862 5186 41914
rect 5198 41862 5250 41914
rect 5262 41862 5314 41914
rect 5326 41862 5378 41914
rect 5390 41862 5442 41914
rect 35854 41862 35906 41914
rect 35918 41862 35970 41914
rect 35982 41862 36034 41914
rect 36046 41862 36098 41914
rect 36110 41862 36162 41914
rect 66574 41862 66626 41914
rect 66638 41862 66690 41914
rect 66702 41862 66754 41914
rect 66766 41862 66818 41914
rect 66830 41862 66882 41914
rect 64880 41760 64932 41812
rect 1216 41556 1268 41608
rect 64604 41599 64656 41608
rect 64604 41565 64613 41599
rect 64613 41565 64647 41599
rect 64647 41565 64656 41599
rect 64604 41556 64656 41565
rect 64788 41599 64840 41608
rect 64788 41565 64797 41599
rect 64797 41565 64831 41599
rect 64831 41565 64840 41599
rect 64788 41556 64840 41565
rect 74356 41599 74408 41608
rect 74356 41565 74365 41599
rect 74365 41565 74399 41599
rect 74399 41565 74408 41599
rect 74356 41556 74408 41565
rect 76380 41599 76432 41608
rect 76380 41565 76389 41599
rect 76389 41565 76423 41599
rect 76423 41565 76432 41599
rect 76380 41556 76432 41565
rect 74632 41531 74684 41540
rect 74632 41497 74641 41531
rect 74641 41497 74675 41531
rect 74675 41497 74684 41531
rect 74632 41488 74684 41497
rect 71228 41463 71280 41472
rect 71228 41429 71237 41463
rect 71237 41429 71271 41463
rect 71271 41429 71280 41463
rect 71228 41420 71280 41429
rect 75920 41420 75972 41472
rect 5794 41318 5846 41370
rect 5858 41318 5910 41370
rect 5922 41318 5974 41370
rect 5986 41318 6038 41370
rect 6050 41318 6102 41370
rect 36514 41318 36566 41370
rect 36578 41318 36630 41370
rect 36642 41318 36694 41370
rect 36706 41318 36758 41370
rect 36770 41318 36822 41370
rect 67234 41318 67286 41370
rect 67298 41318 67350 41370
rect 67362 41318 67414 41370
rect 67426 41318 67478 41370
rect 67490 41318 67542 41370
rect 68284 41080 68336 41132
rect 74356 41216 74408 41268
rect 71228 41148 71280 41200
rect 70492 41055 70544 41064
rect 70492 41021 70501 41055
rect 70501 41021 70535 41055
rect 70535 41021 70544 41055
rect 70492 41012 70544 41021
rect 71136 41012 71188 41064
rect 74632 41012 74684 41064
rect 75920 41055 75972 41064
rect 75920 41021 75929 41055
rect 75929 41021 75963 41055
rect 75963 41021 75972 41055
rect 75920 41012 75972 41021
rect 71964 40919 72016 40928
rect 71964 40885 71973 40919
rect 71973 40885 72007 40919
rect 72007 40885 72016 40919
rect 71964 40876 72016 40885
rect 5134 40774 5186 40826
rect 5198 40774 5250 40826
rect 5262 40774 5314 40826
rect 5326 40774 5378 40826
rect 5390 40774 5442 40826
rect 35854 40774 35906 40826
rect 35918 40774 35970 40826
rect 35982 40774 36034 40826
rect 36046 40774 36098 40826
rect 36110 40774 36162 40826
rect 66574 40774 66626 40826
rect 66638 40774 66690 40826
rect 66702 40774 66754 40826
rect 66766 40774 66818 40826
rect 66830 40774 66882 40826
rect 70492 40672 70544 40724
rect 62672 40604 62724 40656
rect 64788 40604 64840 40656
rect 60924 40579 60976 40588
rect 60924 40545 60933 40579
rect 60933 40545 60967 40579
rect 60967 40545 60976 40579
rect 60924 40536 60976 40545
rect 60832 40511 60884 40520
rect 60832 40477 60841 40511
rect 60841 40477 60875 40511
rect 60875 40477 60884 40511
rect 60832 40468 60884 40477
rect 63500 40536 63552 40588
rect 65156 40536 65208 40588
rect 57612 40400 57664 40452
rect 64788 40468 64840 40520
rect 66168 40536 66220 40588
rect 62120 40400 62172 40452
rect 65984 40511 66036 40520
rect 65984 40477 65993 40511
rect 65993 40477 66027 40511
rect 66027 40477 66036 40511
rect 65984 40468 66036 40477
rect 66076 40511 66128 40520
rect 66076 40477 66085 40511
rect 66085 40477 66119 40511
rect 66119 40477 66128 40511
rect 66076 40468 66128 40477
rect 66904 40604 66956 40656
rect 71504 40604 71556 40656
rect 68284 40579 68336 40588
rect 68284 40545 68293 40579
rect 68293 40545 68327 40579
rect 68327 40545 68336 40579
rect 68284 40536 68336 40545
rect 71136 40579 71188 40588
rect 71136 40545 71145 40579
rect 71145 40545 71179 40579
rect 71179 40545 71188 40579
rect 71136 40536 71188 40545
rect 66996 40400 67048 40452
rect 68008 40443 68060 40452
rect 68008 40409 68017 40443
rect 68017 40409 68051 40443
rect 68051 40409 68060 40443
rect 68008 40400 68060 40409
rect 60924 40332 60976 40384
rect 64604 40332 64656 40384
rect 66444 40332 66496 40384
rect 5794 40230 5846 40282
rect 5858 40230 5910 40282
rect 5922 40230 5974 40282
rect 5986 40230 6038 40282
rect 6050 40230 6102 40282
rect 36514 40230 36566 40282
rect 36578 40230 36630 40282
rect 36642 40230 36694 40282
rect 36706 40230 36758 40282
rect 36770 40230 36822 40282
rect 67234 40230 67286 40282
rect 67298 40230 67350 40282
rect 67362 40230 67414 40282
rect 67426 40230 67478 40282
rect 67490 40230 67542 40282
rect 60832 40128 60884 40180
rect 64604 40128 64656 40180
rect 66076 40128 66128 40180
rect 68008 40128 68060 40180
rect 58992 39992 59044 40044
rect 62120 39992 62172 40044
rect 62672 40035 62724 40044
rect 62672 40001 62681 40035
rect 62681 40001 62715 40035
rect 62715 40001 62724 40035
rect 62672 39992 62724 40001
rect 65984 40035 66036 40044
rect 65984 40001 65993 40035
rect 65993 40001 66027 40035
rect 66027 40001 66036 40035
rect 65984 39992 66036 40001
rect 66168 40103 66220 40112
rect 66168 40069 66177 40103
rect 66177 40069 66211 40103
rect 66211 40069 66220 40103
rect 66168 40060 66220 40069
rect 66904 39992 66956 40044
rect 66996 39992 67048 40044
rect 65800 39788 65852 39840
rect 67088 39924 67140 39976
rect 66444 39856 66496 39908
rect 5134 39686 5186 39738
rect 5198 39686 5250 39738
rect 5262 39686 5314 39738
rect 5326 39686 5378 39738
rect 5390 39686 5442 39738
rect 35854 39686 35906 39738
rect 35918 39686 35970 39738
rect 35982 39686 36034 39738
rect 36046 39686 36098 39738
rect 36110 39686 36162 39738
rect 66574 39686 66626 39738
rect 66638 39686 66690 39738
rect 66702 39686 66754 39738
rect 66766 39686 66818 39738
rect 66830 39686 66882 39738
rect 71136 39584 71188 39636
rect 66168 39516 66220 39568
rect 76196 39559 76248 39568
rect 76196 39525 76205 39559
rect 76205 39525 76239 39559
rect 76239 39525 76248 39559
rect 76196 39516 76248 39525
rect 57612 39448 57664 39500
rect 58348 39380 58400 39432
rect 58992 39380 59044 39432
rect 66260 39380 66312 39432
rect 66904 39380 66956 39432
rect 75736 39380 75788 39432
rect 57060 39355 57112 39364
rect 57060 39321 57069 39355
rect 57069 39321 57103 39355
rect 57103 39321 57112 39355
rect 57060 39312 57112 39321
rect 70676 39312 70728 39364
rect 71596 39312 71648 39364
rect 75828 39312 75880 39364
rect 57980 39244 58032 39296
rect 66904 39287 66956 39296
rect 66904 39253 66913 39287
rect 66913 39253 66947 39287
rect 66947 39253 66956 39287
rect 66904 39244 66956 39253
rect 67088 39287 67140 39296
rect 67088 39253 67097 39287
rect 67097 39253 67131 39287
rect 67131 39253 67140 39287
rect 67088 39244 67140 39253
rect 71044 39287 71096 39296
rect 71044 39253 71053 39287
rect 71053 39253 71087 39287
rect 71087 39253 71096 39287
rect 71044 39244 71096 39253
rect 71228 39287 71280 39296
rect 71228 39253 71237 39287
rect 71237 39253 71271 39287
rect 71271 39253 71280 39287
rect 71228 39244 71280 39253
rect 76012 39287 76064 39296
rect 76012 39253 76021 39287
rect 76021 39253 76055 39287
rect 76055 39253 76064 39287
rect 76012 39244 76064 39253
rect 5794 39142 5846 39194
rect 5858 39142 5910 39194
rect 5922 39142 5974 39194
rect 5986 39142 6038 39194
rect 6050 39142 6102 39194
rect 36514 39142 36566 39194
rect 36578 39142 36630 39194
rect 36642 39142 36694 39194
rect 36706 39142 36758 39194
rect 36770 39142 36822 39194
rect 67234 39142 67286 39194
rect 67298 39142 67350 39194
rect 67362 39142 67414 39194
rect 67426 39142 67478 39194
rect 67490 39142 67542 39194
rect 71136 39083 71188 39092
rect 71136 39049 71145 39083
rect 71145 39049 71179 39083
rect 71179 39049 71188 39083
rect 71136 39040 71188 39049
rect 71504 39083 71556 39092
rect 71504 39049 71513 39083
rect 71513 39049 71547 39083
rect 71547 39049 71556 39083
rect 71504 39040 71556 39049
rect 71596 39083 71648 39092
rect 71596 39049 71605 39083
rect 71605 39049 71639 39083
rect 71639 39049 71648 39083
rect 71596 39040 71648 39049
rect 75920 39040 75972 39092
rect 1308 38904 1360 38956
rect 71044 38904 71096 38956
rect 71964 38947 72016 38956
rect 71964 38913 71973 38947
rect 71973 38913 72007 38947
rect 72007 38913 72016 38947
rect 71964 38904 72016 38913
rect 74632 38904 74684 38956
rect 70676 38836 70728 38888
rect 76288 38904 76340 38956
rect 75736 38836 75788 38888
rect 77484 38811 77536 38820
rect 77484 38777 77493 38811
rect 77493 38777 77527 38811
rect 77527 38777 77536 38811
rect 77484 38768 77536 38777
rect 66444 38700 66496 38752
rect 75368 38700 75420 38752
rect 75828 38700 75880 38752
rect 5134 38598 5186 38650
rect 5198 38598 5250 38650
rect 5262 38598 5314 38650
rect 5326 38598 5378 38650
rect 5390 38598 5442 38650
rect 35854 38598 35906 38650
rect 35918 38598 35970 38650
rect 35982 38598 36034 38650
rect 36046 38598 36098 38650
rect 36110 38598 36162 38650
rect 66574 38598 66626 38650
rect 66638 38598 66690 38650
rect 66702 38598 66754 38650
rect 66766 38598 66818 38650
rect 66830 38598 66882 38650
rect 57060 38539 57112 38548
rect 57060 38505 57069 38539
rect 57069 38505 57103 38539
rect 57103 38505 57112 38539
rect 57060 38496 57112 38505
rect 63500 38496 63552 38548
rect 68284 38496 68336 38548
rect 68928 38496 68980 38548
rect 76012 38496 76064 38548
rect 76288 38539 76340 38548
rect 76288 38505 76297 38539
rect 76297 38505 76331 38539
rect 76331 38505 76340 38539
rect 76288 38496 76340 38505
rect 57336 38335 57388 38344
rect 57336 38301 57345 38335
rect 57345 38301 57379 38335
rect 57379 38301 57388 38335
rect 57336 38292 57388 38301
rect 74632 38335 74684 38344
rect 74632 38301 74641 38335
rect 74641 38301 74675 38335
rect 74675 38301 74684 38335
rect 74632 38292 74684 38301
rect 76104 38335 76156 38344
rect 76104 38301 76113 38335
rect 76113 38301 76147 38335
rect 76147 38301 76156 38335
rect 76104 38292 76156 38301
rect 76288 38292 76340 38344
rect 57796 38267 57848 38276
rect 57796 38233 57805 38267
rect 57805 38233 57839 38267
rect 57839 38233 57848 38267
rect 57796 38224 57848 38233
rect 57980 38267 58032 38276
rect 57980 38233 57989 38267
rect 57989 38233 58023 38267
rect 58023 38233 58032 38267
rect 57980 38224 58032 38233
rect 66444 38224 66496 38276
rect 77484 38199 77536 38208
rect 77484 38165 77493 38199
rect 77493 38165 77527 38199
rect 77527 38165 77536 38199
rect 77484 38156 77536 38165
rect 5794 38054 5846 38106
rect 5858 38054 5910 38106
rect 5922 38054 5974 38106
rect 5986 38054 6038 38106
rect 6050 38054 6102 38106
rect 36514 38054 36566 38106
rect 36578 38054 36630 38106
rect 36642 38054 36694 38106
rect 36706 38054 36758 38106
rect 36770 38054 36822 38106
rect 67234 38054 67286 38106
rect 67298 38054 67350 38106
rect 67362 38054 67414 38106
rect 67426 38054 67478 38106
rect 67490 38054 67542 38106
rect 68284 37884 68336 37936
rect 76472 37816 76524 37868
rect 77484 37655 77536 37664
rect 77484 37621 77493 37655
rect 77493 37621 77527 37655
rect 77527 37621 77536 37655
rect 77484 37612 77536 37621
rect 5134 37510 5186 37562
rect 5198 37510 5250 37562
rect 5262 37510 5314 37562
rect 5326 37510 5378 37562
rect 5390 37510 5442 37562
rect 35854 37510 35906 37562
rect 35918 37510 35970 37562
rect 35982 37510 36034 37562
rect 36046 37510 36098 37562
rect 36110 37510 36162 37562
rect 66574 37510 66626 37562
rect 66638 37510 66690 37562
rect 66702 37510 66754 37562
rect 66766 37510 66818 37562
rect 66830 37510 66882 37562
rect 63500 37272 63552 37324
rect 65340 37272 65392 37324
rect 57796 37204 57848 37256
rect 60004 37204 60056 37256
rect 66904 37204 66956 37256
rect 75368 37247 75420 37256
rect 75368 37213 75377 37247
rect 75377 37213 75411 37247
rect 75411 37213 75420 37247
rect 75368 37204 75420 37213
rect 57980 37136 58032 37188
rect 65984 37136 66036 37188
rect 56784 37068 56836 37120
rect 57336 37068 57388 37120
rect 76104 37136 76156 37188
rect 66536 37111 66588 37120
rect 66536 37077 66545 37111
rect 66545 37077 66579 37111
rect 66579 37077 66588 37111
rect 66536 37068 66588 37077
rect 77484 37111 77536 37120
rect 77484 37077 77493 37111
rect 77493 37077 77527 37111
rect 77527 37077 77536 37111
rect 77484 37068 77536 37077
rect 5794 36966 5846 37018
rect 5858 36966 5910 37018
rect 5922 36966 5974 37018
rect 5986 36966 6038 37018
rect 6050 36966 6102 37018
rect 36514 36966 36566 37018
rect 36578 36966 36630 37018
rect 36642 36966 36694 37018
rect 36706 36966 36758 37018
rect 36770 36966 36822 37018
rect 67234 36966 67286 37018
rect 67298 36966 67350 37018
rect 67362 36966 67414 37018
rect 67426 36966 67478 37018
rect 67490 36966 67542 37018
rect 65340 36864 65392 36916
rect 65984 36864 66036 36916
rect 60004 36839 60056 36848
rect 60004 36805 60013 36839
rect 60013 36805 60047 36839
rect 60047 36805 60056 36839
rect 60004 36796 60056 36805
rect 60372 36839 60424 36848
rect 60372 36805 60381 36839
rect 60381 36805 60415 36839
rect 60415 36805 60424 36839
rect 60372 36796 60424 36805
rect 60924 36796 60976 36848
rect 57980 36728 58032 36780
rect 60188 36771 60240 36780
rect 60188 36737 60197 36771
rect 60197 36737 60231 36771
rect 60231 36737 60240 36771
rect 60188 36728 60240 36737
rect 60280 36771 60332 36780
rect 60280 36737 60289 36771
rect 60289 36737 60323 36771
rect 60323 36737 60332 36771
rect 60280 36728 60332 36737
rect 65616 36771 65668 36780
rect 65616 36737 65625 36771
rect 65625 36737 65659 36771
rect 65659 36737 65668 36771
rect 65616 36728 65668 36737
rect 65800 36771 65852 36780
rect 65800 36737 65809 36771
rect 65809 36737 65843 36771
rect 65843 36737 65852 36771
rect 65800 36728 65852 36737
rect 66536 36796 66588 36848
rect 66168 36771 66220 36780
rect 66168 36737 66177 36771
rect 66177 36737 66211 36771
rect 66211 36737 66220 36771
rect 66168 36728 66220 36737
rect 66996 36728 67048 36780
rect 5134 36422 5186 36474
rect 5198 36422 5250 36474
rect 5262 36422 5314 36474
rect 5326 36422 5378 36474
rect 5390 36422 5442 36474
rect 35854 36422 35906 36474
rect 35918 36422 35970 36474
rect 35982 36422 36034 36474
rect 36046 36422 36098 36474
rect 36110 36422 36162 36474
rect 66574 36422 66626 36474
rect 66638 36422 66690 36474
rect 66702 36422 66754 36474
rect 66766 36422 66818 36474
rect 66830 36422 66882 36474
rect 65616 36320 65668 36372
rect 65984 36320 66036 36372
rect 76472 36363 76524 36372
rect 76472 36329 76481 36363
rect 76481 36329 76515 36363
rect 76515 36329 76524 36363
rect 76472 36320 76524 36329
rect 60004 36252 60056 36304
rect 60188 36227 60240 36236
rect 60188 36193 60197 36227
rect 60197 36193 60231 36227
rect 60231 36193 60240 36227
rect 60188 36184 60240 36193
rect 60280 36227 60332 36236
rect 60280 36193 60289 36227
rect 60289 36193 60323 36227
rect 60323 36193 60332 36227
rect 60280 36184 60332 36193
rect 60924 36184 60976 36236
rect 67088 36116 67140 36168
rect 71688 36184 71740 36236
rect 76380 36184 76432 36236
rect 60372 36048 60424 36100
rect 70676 36091 70728 36100
rect 60556 36023 60608 36032
rect 60556 35989 60565 36023
rect 60565 35989 60599 36023
rect 60599 35989 60608 36023
rect 60556 35980 60608 35989
rect 70676 36057 70685 36091
rect 70685 36057 70719 36091
rect 70719 36057 70728 36091
rect 70676 36048 70728 36057
rect 70860 36159 70912 36168
rect 70860 36125 70869 36159
rect 70869 36125 70903 36159
rect 70903 36125 70912 36159
rect 70860 36116 70912 36125
rect 71044 36116 71096 36168
rect 73160 36116 73212 36168
rect 74080 36159 74132 36168
rect 74080 36125 74089 36159
rect 74089 36125 74123 36159
rect 74123 36125 74132 36159
rect 74080 36116 74132 36125
rect 76196 36159 76248 36168
rect 76196 36125 76205 36159
rect 76205 36125 76239 36159
rect 76239 36125 76248 36159
rect 76196 36116 76248 36125
rect 76288 36159 76340 36168
rect 76288 36125 76297 36159
rect 76297 36125 76331 36159
rect 76331 36125 76340 36159
rect 76288 36116 76340 36125
rect 71136 36048 71188 36100
rect 62120 35980 62172 36032
rect 75828 36023 75880 36032
rect 75828 35989 75837 36023
rect 75837 35989 75871 36023
rect 75871 35989 75880 36023
rect 75828 35980 75880 35989
rect 5794 35878 5846 35930
rect 5858 35878 5910 35930
rect 5922 35878 5974 35930
rect 5986 35878 6038 35930
rect 6050 35878 6102 35930
rect 36514 35878 36566 35930
rect 36578 35878 36630 35930
rect 36642 35878 36694 35930
rect 36706 35878 36758 35930
rect 36770 35878 36822 35930
rect 67234 35878 67286 35930
rect 67298 35878 67350 35930
rect 67362 35878 67414 35930
rect 67426 35878 67478 35930
rect 67490 35878 67542 35930
rect 58072 35683 58124 35692
rect 58072 35649 58081 35683
rect 58081 35649 58115 35683
rect 58115 35649 58124 35683
rect 58072 35640 58124 35649
rect 60280 35640 60332 35692
rect 63500 35776 63552 35828
rect 73160 35776 73212 35828
rect 60556 35708 60608 35760
rect 70676 35708 70728 35760
rect 56784 35615 56836 35624
rect 56784 35581 56793 35615
rect 56793 35581 56827 35615
rect 56827 35581 56836 35615
rect 56784 35572 56836 35581
rect 60372 35615 60424 35624
rect 60372 35581 60381 35615
rect 60381 35581 60415 35615
rect 60415 35581 60424 35615
rect 60372 35572 60424 35581
rect 66168 35640 66220 35692
rect 71136 35683 71188 35692
rect 71136 35649 71145 35683
rect 71145 35649 71179 35683
rect 71179 35649 71188 35683
rect 71136 35640 71188 35649
rect 71688 35683 71740 35692
rect 71688 35649 71697 35683
rect 71697 35649 71731 35683
rect 71731 35649 71740 35683
rect 71688 35640 71740 35649
rect 75828 35640 75880 35692
rect 58348 35504 58400 35556
rect 62120 35615 62172 35624
rect 62120 35581 62129 35615
rect 62129 35581 62163 35615
rect 62163 35581 62172 35615
rect 62120 35572 62172 35581
rect 70124 35615 70176 35624
rect 70124 35581 70133 35615
rect 70133 35581 70167 35615
rect 70167 35581 70176 35615
rect 70124 35572 70176 35581
rect 70676 35504 70728 35556
rect 1216 35436 1268 35488
rect 56416 35479 56468 35488
rect 56416 35445 56425 35479
rect 56425 35445 56459 35479
rect 56459 35445 56468 35479
rect 56416 35436 56468 35445
rect 71320 35436 71372 35488
rect 5134 35334 5186 35386
rect 5198 35334 5250 35386
rect 5262 35334 5314 35386
rect 5326 35334 5378 35386
rect 5390 35334 5442 35386
rect 35854 35334 35906 35386
rect 35918 35334 35970 35386
rect 35982 35334 36034 35386
rect 36046 35334 36098 35386
rect 36110 35334 36162 35386
rect 66574 35334 66626 35386
rect 66638 35334 66690 35386
rect 66702 35334 66754 35386
rect 66766 35334 66818 35386
rect 66830 35334 66882 35386
rect 56416 35232 56468 35284
rect 58072 35275 58124 35284
rect 58072 35241 58081 35275
rect 58081 35241 58115 35275
rect 58115 35241 58124 35275
rect 58072 35232 58124 35241
rect 70860 35232 70912 35284
rect 60372 35096 60424 35148
rect 70124 35096 70176 35148
rect 58348 35071 58400 35080
rect 58348 35037 58357 35071
rect 58357 35037 58391 35071
rect 58391 35037 58400 35071
rect 58348 35028 58400 35037
rect 66996 35028 67048 35080
rect 70676 35071 70728 35080
rect 70676 35037 70685 35071
rect 70685 35037 70719 35071
rect 70719 35037 70728 35071
rect 70676 35028 70728 35037
rect 5794 34790 5846 34842
rect 5858 34790 5910 34842
rect 5922 34790 5974 34842
rect 5986 34790 6038 34842
rect 6050 34790 6102 34842
rect 36514 34790 36566 34842
rect 36578 34790 36630 34842
rect 36642 34790 36694 34842
rect 36706 34790 36758 34842
rect 36770 34790 36822 34842
rect 67234 34790 67286 34842
rect 67298 34790 67350 34842
rect 67362 34790 67414 34842
rect 67426 34790 67478 34842
rect 67490 34790 67542 34842
rect 68928 34688 68980 34740
rect 70308 34620 70360 34672
rect 71320 34663 71372 34672
rect 71320 34629 71329 34663
rect 71329 34629 71363 34663
rect 71363 34629 71372 34663
rect 71320 34620 71372 34629
rect 66996 34595 67048 34604
rect 66996 34561 67005 34595
rect 67005 34561 67039 34595
rect 67039 34561 67048 34595
rect 66996 34552 67048 34561
rect 74080 34620 74132 34672
rect 76196 34620 76248 34672
rect 77484 34595 77536 34604
rect 77484 34561 77493 34595
rect 77493 34561 77527 34595
rect 77527 34561 77536 34595
rect 77484 34552 77536 34561
rect 65984 34527 66036 34536
rect 65984 34493 65993 34527
rect 65993 34493 66027 34527
rect 66027 34493 66036 34527
rect 65984 34484 66036 34493
rect 70124 34484 70176 34536
rect 71872 34527 71924 34536
rect 71872 34493 71881 34527
rect 71881 34493 71915 34527
rect 71915 34493 71924 34527
rect 71872 34484 71924 34493
rect 68008 34348 68060 34400
rect 5134 34246 5186 34298
rect 5198 34246 5250 34298
rect 5262 34246 5314 34298
rect 5326 34246 5378 34298
rect 5390 34246 5442 34298
rect 35854 34246 35906 34298
rect 35918 34246 35970 34298
rect 35982 34246 36034 34298
rect 36046 34246 36098 34298
rect 36110 34246 36162 34298
rect 66574 34246 66626 34298
rect 66638 34246 66690 34298
rect 66702 34246 66754 34298
rect 66766 34246 66818 34298
rect 66830 34246 66882 34298
rect 66996 34144 67048 34196
rect 70308 34144 70360 34196
rect 68008 34051 68060 34060
rect 68008 34017 68017 34051
rect 68017 34017 68051 34051
rect 68051 34017 68060 34051
rect 68008 34008 68060 34017
rect 68928 34008 68980 34060
rect 66904 33940 66956 33992
rect 66260 33804 66312 33856
rect 71872 33940 71924 33992
rect 5794 33702 5846 33754
rect 5858 33702 5910 33754
rect 5922 33702 5974 33754
rect 5986 33702 6038 33754
rect 6050 33702 6102 33754
rect 36514 33702 36566 33754
rect 36578 33702 36630 33754
rect 36642 33702 36694 33754
rect 36706 33702 36758 33754
rect 36770 33702 36822 33754
rect 67234 33702 67286 33754
rect 67298 33702 67350 33754
rect 67362 33702 67414 33754
rect 67426 33702 67478 33754
rect 67490 33702 67542 33754
rect 66904 33643 66956 33652
rect 66904 33609 66913 33643
rect 66913 33609 66947 33643
rect 66947 33609 66956 33643
rect 66904 33600 66956 33609
rect 66260 33464 66312 33516
rect 5134 33158 5186 33210
rect 5198 33158 5250 33210
rect 5262 33158 5314 33210
rect 5326 33158 5378 33210
rect 5390 33158 5442 33210
rect 35854 33158 35906 33210
rect 35918 33158 35970 33210
rect 35982 33158 36034 33210
rect 36046 33158 36098 33210
rect 36110 33158 36162 33210
rect 66574 33158 66626 33210
rect 66638 33158 66690 33210
rect 66702 33158 66754 33210
rect 66766 33158 66818 33210
rect 66830 33158 66882 33210
rect 5794 32614 5846 32666
rect 5858 32614 5910 32666
rect 5922 32614 5974 32666
rect 5986 32614 6038 32666
rect 6050 32614 6102 32666
rect 36514 32614 36566 32666
rect 36578 32614 36630 32666
rect 36642 32614 36694 32666
rect 36706 32614 36758 32666
rect 36770 32614 36822 32666
rect 67234 32614 67286 32666
rect 67298 32614 67350 32666
rect 67362 32614 67414 32666
rect 67426 32614 67478 32666
rect 67490 32614 67542 32666
rect 1216 32172 1268 32224
rect 5134 32070 5186 32122
rect 5198 32070 5250 32122
rect 5262 32070 5314 32122
rect 5326 32070 5378 32122
rect 5390 32070 5442 32122
rect 35854 32070 35906 32122
rect 35918 32070 35970 32122
rect 35982 32070 36034 32122
rect 36046 32070 36098 32122
rect 36110 32070 36162 32122
rect 66574 32070 66626 32122
rect 66638 32070 66690 32122
rect 66702 32070 66754 32122
rect 66766 32070 66818 32122
rect 66830 32070 66882 32122
rect 5794 31526 5846 31578
rect 5858 31526 5910 31578
rect 5922 31526 5974 31578
rect 5986 31526 6038 31578
rect 6050 31526 6102 31578
rect 36514 31526 36566 31578
rect 36578 31526 36630 31578
rect 36642 31526 36694 31578
rect 36706 31526 36758 31578
rect 36770 31526 36822 31578
rect 67234 31526 67286 31578
rect 67298 31526 67350 31578
rect 67362 31526 67414 31578
rect 67426 31526 67478 31578
rect 67490 31526 67542 31578
rect 5134 30982 5186 31034
rect 5198 30982 5250 31034
rect 5262 30982 5314 31034
rect 5326 30982 5378 31034
rect 5390 30982 5442 31034
rect 35854 30982 35906 31034
rect 35918 30982 35970 31034
rect 35982 30982 36034 31034
rect 36046 30982 36098 31034
rect 36110 30982 36162 31034
rect 66574 30982 66626 31034
rect 66638 30982 66690 31034
rect 66702 30982 66754 31034
rect 66766 30982 66818 31034
rect 66830 30982 66882 31034
rect 5794 30438 5846 30490
rect 5858 30438 5910 30490
rect 5922 30438 5974 30490
rect 5986 30438 6038 30490
rect 6050 30438 6102 30490
rect 36514 30438 36566 30490
rect 36578 30438 36630 30490
rect 36642 30438 36694 30490
rect 36706 30438 36758 30490
rect 36770 30438 36822 30490
rect 67234 30438 67286 30490
rect 67298 30438 67350 30490
rect 67362 30438 67414 30490
rect 67426 30438 67478 30490
rect 67490 30438 67542 30490
rect 5134 29894 5186 29946
rect 5198 29894 5250 29946
rect 5262 29894 5314 29946
rect 5326 29894 5378 29946
rect 5390 29894 5442 29946
rect 35854 29894 35906 29946
rect 35918 29894 35970 29946
rect 35982 29894 36034 29946
rect 36046 29894 36098 29946
rect 36110 29894 36162 29946
rect 66574 29894 66626 29946
rect 66638 29894 66690 29946
rect 66702 29894 66754 29946
rect 66766 29894 66818 29946
rect 66830 29894 66882 29946
rect 5794 29350 5846 29402
rect 5858 29350 5910 29402
rect 5922 29350 5974 29402
rect 5986 29350 6038 29402
rect 6050 29350 6102 29402
rect 36514 29350 36566 29402
rect 36578 29350 36630 29402
rect 36642 29350 36694 29402
rect 36706 29350 36758 29402
rect 36770 29350 36822 29402
rect 67234 29350 67286 29402
rect 67298 29350 67350 29402
rect 67362 29350 67414 29402
rect 67426 29350 67478 29402
rect 67490 29350 67542 29402
rect 2320 29019 2372 29028
rect 2320 28985 2329 29019
rect 2329 28985 2363 29019
rect 2363 28985 2372 29019
rect 2320 28976 2372 28985
rect 5134 28806 5186 28858
rect 5198 28806 5250 28858
rect 5262 28806 5314 28858
rect 5326 28806 5378 28858
rect 5390 28806 5442 28858
rect 35854 28806 35906 28858
rect 35918 28806 35970 28858
rect 35982 28806 36034 28858
rect 36046 28806 36098 28858
rect 36110 28806 36162 28858
rect 66574 28806 66626 28858
rect 66638 28806 66690 28858
rect 66702 28806 66754 28858
rect 66766 28806 66818 28858
rect 66830 28806 66882 28858
rect 5794 28262 5846 28314
rect 5858 28262 5910 28314
rect 5922 28262 5974 28314
rect 5986 28262 6038 28314
rect 6050 28262 6102 28314
rect 36514 28262 36566 28314
rect 36578 28262 36630 28314
rect 36642 28262 36694 28314
rect 36706 28262 36758 28314
rect 36770 28262 36822 28314
rect 67234 28262 67286 28314
rect 67298 28262 67350 28314
rect 67362 28262 67414 28314
rect 67426 28262 67478 28314
rect 67490 28262 67542 28314
rect 1216 27956 1268 28008
rect 5134 27718 5186 27770
rect 5198 27718 5250 27770
rect 5262 27718 5314 27770
rect 5326 27718 5378 27770
rect 5390 27718 5442 27770
rect 35854 27718 35906 27770
rect 35918 27718 35970 27770
rect 35982 27718 36034 27770
rect 36046 27718 36098 27770
rect 36110 27718 36162 27770
rect 66574 27718 66626 27770
rect 66638 27718 66690 27770
rect 66702 27718 66754 27770
rect 66766 27718 66818 27770
rect 66830 27718 66882 27770
rect 5794 27174 5846 27226
rect 5858 27174 5910 27226
rect 5922 27174 5974 27226
rect 5986 27174 6038 27226
rect 6050 27174 6102 27226
rect 36514 27174 36566 27226
rect 36578 27174 36630 27226
rect 36642 27174 36694 27226
rect 36706 27174 36758 27226
rect 36770 27174 36822 27226
rect 67234 27174 67286 27226
rect 67298 27174 67350 27226
rect 67362 27174 67414 27226
rect 67426 27174 67478 27226
rect 67490 27174 67542 27226
rect 1216 26732 1268 26784
rect 5134 26630 5186 26682
rect 5198 26630 5250 26682
rect 5262 26630 5314 26682
rect 5326 26630 5378 26682
rect 5390 26630 5442 26682
rect 35854 26630 35906 26682
rect 35918 26630 35970 26682
rect 35982 26630 36034 26682
rect 36046 26630 36098 26682
rect 36110 26630 36162 26682
rect 66574 26630 66626 26682
rect 66638 26630 66690 26682
rect 66702 26630 66754 26682
rect 66766 26630 66818 26682
rect 66830 26630 66882 26682
rect 2320 26367 2372 26376
rect 2320 26333 2329 26367
rect 2329 26333 2363 26367
rect 2363 26333 2372 26367
rect 2320 26324 2372 26333
rect 5794 26086 5846 26138
rect 5858 26086 5910 26138
rect 5922 26086 5974 26138
rect 5986 26086 6038 26138
rect 6050 26086 6102 26138
rect 36514 26086 36566 26138
rect 36578 26086 36630 26138
rect 36642 26086 36694 26138
rect 36706 26086 36758 26138
rect 36770 26086 36822 26138
rect 67234 26086 67286 26138
rect 67298 26086 67350 26138
rect 67362 26086 67414 26138
rect 67426 26086 67478 26138
rect 67490 26086 67542 26138
rect 5134 25542 5186 25594
rect 5198 25542 5250 25594
rect 5262 25542 5314 25594
rect 5326 25542 5378 25594
rect 5390 25542 5442 25594
rect 35854 25542 35906 25594
rect 35918 25542 35970 25594
rect 35982 25542 36034 25594
rect 36046 25542 36098 25594
rect 36110 25542 36162 25594
rect 66574 25542 66626 25594
rect 66638 25542 66690 25594
rect 66702 25542 66754 25594
rect 66766 25542 66818 25594
rect 66830 25542 66882 25594
rect 5794 24998 5846 25050
rect 5858 24998 5910 25050
rect 5922 24998 5974 25050
rect 5986 24998 6038 25050
rect 6050 24998 6102 25050
rect 36514 24998 36566 25050
rect 36578 24998 36630 25050
rect 36642 24998 36694 25050
rect 36706 24998 36758 25050
rect 36770 24998 36822 25050
rect 67234 24998 67286 25050
rect 67298 24998 67350 25050
rect 67362 24998 67414 25050
rect 67426 24998 67478 25050
rect 67490 24998 67542 25050
rect 5134 24454 5186 24506
rect 5198 24454 5250 24506
rect 5262 24454 5314 24506
rect 5326 24454 5378 24506
rect 5390 24454 5442 24506
rect 35854 24454 35906 24506
rect 35918 24454 35970 24506
rect 35982 24454 36034 24506
rect 36046 24454 36098 24506
rect 36110 24454 36162 24506
rect 66574 24454 66626 24506
rect 66638 24454 66690 24506
rect 66702 24454 66754 24506
rect 66766 24454 66818 24506
rect 66830 24454 66882 24506
rect 5794 23910 5846 23962
rect 5858 23910 5910 23962
rect 5922 23910 5974 23962
rect 5986 23910 6038 23962
rect 6050 23910 6102 23962
rect 36514 23910 36566 23962
rect 36578 23910 36630 23962
rect 36642 23910 36694 23962
rect 36706 23910 36758 23962
rect 36770 23910 36822 23962
rect 67234 23910 67286 23962
rect 67298 23910 67350 23962
rect 67362 23910 67414 23962
rect 67426 23910 67478 23962
rect 67490 23910 67542 23962
rect 2320 23511 2372 23520
rect 2320 23477 2329 23511
rect 2329 23477 2363 23511
rect 2363 23477 2372 23511
rect 2320 23468 2372 23477
rect 5134 23366 5186 23418
rect 5198 23366 5250 23418
rect 5262 23366 5314 23418
rect 5326 23366 5378 23418
rect 5390 23366 5442 23418
rect 35854 23366 35906 23418
rect 35918 23366 35970 23418
rect 35982 23366 36034 23418
rect 36046 23366 36098 23418
rect 36110 23366 36162 23418
rect 66574 23366 66626 23418
rect 66638 23366 66690 23418
rect 66702 23366 66754 23418
rect 66766 23366 66818 23418
rect 66830 23366 66882 23418
rect 5794 22822 5846 22874
rect 5858 22822 5910 22874
rect 5922 22822 5974 22874
rect 5986 22822 6038 22874
rect 6050 22822 6102 22874
rect 36514 22822 36566 22874
rect 36578 22822 36630 22874
rect 36642 22822 36694 22874
rect 36706 22822 36758 22874
rect 36770 22822 36822 22874
rect 67234 22822 67286 22874
rect 67298 22822 67350 22874
rect 67362 22822 67414 22874
rect 67426 22822 67478 22874
rect 67490 22822 67542 22874
rect 5134 22278 5186 22330
rect 5198 22278 5250 22330
rect 5262 22278 5314 22330
rect 5326 22278 5378 22330
rect 5390 22278 5442 22330
rect 35854 22278 35906 22330
rect 35918 22278 35970 22330
rect 35982 22278 36034 22330
rect 36046 22278 36098 22330
rect 36110 22278 36162 22330
rect 66574 22278 66626 22330
rect 66638 22278 66690 22330
rect 66702 22278 66754 22330
rect 66766 22278 66818 22330
rect 66830 22278 66882 22330
rect 5794 21734 5846 21786
rect 5858 21734 5910 21786
rect 5922 21734 5974 21786
rect 5986 21734 6038 21786
rect 6050 21734 6102 21786
rect 36514 21734 36566 21786
rect 36578 21734 36630 21786
rect 36642 21734 36694 21786
rect 36706 21734 36758 21786
rect 36770 21734 36822 21786
rect 67234 21734 67286 21786
rect 67298 21734 67350 21786
rect 67362 21734 67414 21786
rect 67426 21734 67478 21786
rect 67490 21734 67542 21786
rect 77576 21335 77628 21344
rect 77576 21301 77585 21335
rect 77585 21301 77619 21335
rect 77619 21301 77628 21335
rect 77576 21292 77628 21301
rect 5134 21190 5186 21242
rect 5198 21190 5250 21242
rect 5262 21190 5314 21242
rect 5326 21190 5378 21242
rect 5390 21190 5442 21242
rect 35854 21190 35906 21242
rect 35918 21190 35970 21242
rect 35982 21190 36034 21242
rect 36046 21190 36098 21242
rect 36110 21190 36162 21242
rect 66574 21190 66626 21242
rect 66638 21190 66690 21242
rect 66702 21190 66754 21242
rect 66766 21190 66818 21242
rect 66830 21190 66882 21242
rect 5794 20646 5846 20698
rect 5858 20646 5910 20698
rect 5922 20646 5974 20698
rect 5986 20646 6038 20698
rect 6050 20646 6102 20698
rect 36514 20646 36566 20698
rect 36578 20646 36630 20698
rect 36642 20646 36694 20698
rect 36706 20646 36758 20698
rect 36770 20646 36822 20698
rect 67234 20646 67286 20698
rect 67298 20646 67350 20698
rect 67362 20646 67414 20698
rect 67426 20646 67478 20698
rect 67490 20646 67542 20698
rect 5134 20102 5186 20154
rect 5198 20102 5250 20154
rect 5262 20102 5314 20154
rect 5326 20102 5378 20154
rect 5390 20102 5442 20154
rect 35854 20102 35906 20154
rect 35918 20102 35970 20154
rect 35982 20102 36034 20154
rect 36046 20102 36098 20154
rect 36110 20102 36162 20154
rect 66574 20102 66626 20154
rect 66638 20102 66690 20154
rect 66702 20102 66754 20154
rect 66766 20102 66818 20154
rect 66830 20102 66882 20154
rect 5794 19558 5846 19610
rect 5858 19558 5910 19610
rect 5922 19558 5974 19610
rect 5986 19558 6038 19610
rect 6050 19558 6102 19610
rect 36514 19558 36566 19610
rect 36578 19558 36630 19610
rect 36642 19558 36694 19610
rect 36706 19558 36758 19610
rect 36770 19558 36822 19610
rect 67234 19558 67286 19610
rect 67298 19558 67350 19610
rect 67362 19558 67414 19610
rect 67426 19558 67478 19610
rect 67490 19558 67542 19610
rect 5134 19014 5186 19066
rect 5198 19014 5250 19066
rect 5262 19014 5314 19066
rect 5326 19014 5378 19066
rect 5390 19014 5442 19066
rect 35854 19014 35906 19066
rect 35918 19014 35970 19066
rect 35982 19014 36034 19066
rect 36046 19014 36098 19066
rect 36110 19014 36162 19066
rect 66574 19014 66626 19066
rect 66638 19014 66690 19066
rect 66702 19014 66754 19066
rect 66766 19014 66818 19066
rect 66830 19014 66882 19066
rect 5794 18470 5846 18522
rect 5858 18470 5910 18522
rect 5922 18470 5974 18522
rect 5986 18470 6038 18522
rect 6050 18470 6102 18522
rect 36514 18470 36566 18522
rect 36578 18470 36630 18522
rect 36642 18470 36694 18522
rect 36706 18470 36758 18522
rect 36770 18470 36822 18522
rect 67234 18470 67286 18522
rect 67298 18470 67350 18522
rect 67362 18470 67414 18522
rect 67426 18470 67478 18522
rect 67490 18470 67542 18522
rect 5134 17926 5186 17978
rect 5198 17926 5250 17978
rect 5262 17926 5314 17978
rect 5326 17926 5378 17978
rect 5390 17926 5442 17978
rect 35854 17926 35906 17978
rect 35918 17926 35970 17978
rect 35982 17926 36034 17978
rect 36046 17926 36098 17978
rect 36110 17926 36162 17978
rect 66574 17926 66626 17978
rect 66638 17926 66690 17978
rect 66702 17926 66754 17978
rect 66766 17926 66818 17978
rect 66830 17926 66882 17978
rect 5794 17382 5846 17434
rect 5858 17382 5910 17434
rect 5922 17382 5974 17434
rect 5986 17382 6038 17434
rect 6050 17382 6102 17434
rect 36514 17382 36566 17434
rect 36578 17382 36630 17434
rect 36642 17382 36694 17434
rect 36706 17382 36758 17434
rect 36770 17382 36822 17434
rect 67234 17382 67286 17434
rect 67298 17382 67350 17434
rect 67362 17382 67414 17434
rect 67426 17382 67478 17434
rect 67490 17382 67542 17434
rect 5134 16838 5186 16890
rect 5198 16838 5250 16890
rect 5262 16838 5314 16890
rect 5326 16838 5378 16890
rect 5390 16838 5442 16890
rect 35854 16838 35906 16890
rect 35918 16838 35970 16890
rect 35982 16838 36034 16890
rect 36046 16838 36098 16890
rect 36110 16838 36162 16890
rect 66574 16838 66626 16890
rect 66638 16838 66690 16890
rect 66702 16838 66754 16890
rect 66766 16838 66818 16890
rect 66830 16838 66882 16890
rect 77576 16643 77628 16652
rect 77576 16609 77585 16643
rect 77585 16609 77619 16643
rect 77619 16609 77628 16643
rect 77576 16600 77628 16609
rect 5794 16294 5846 16346
rect 5858 16294 5910 16346
rect 5922 16294 5974 16346
rect 5986 16294 6038 16346
rect 6050 16294 6102 16346
rect 36514 16294 36566 16346
rect 36578 16294 36630 16346
rect 36642 16294 36694 16346
rect 36706 16294 36758 16346
rect 36770 16294 36822 16346
rect 67234 16294 67286 16346
rect 67298 16294 67350 16346
rect 67362 16294 67414 16346
rect 67426 16294 67478 16346
rect 67490 16294 67542 16346
rect 5134 15750 5186 15802
rect 5198 15750 5250 15802
rect 5262 15750 5314 15802
rect 5326 15750 5378 15802
rect 5390 15750 5442 15802
rect 35854 15750 35906 15802
rect 35918 15750 35970 15802
rect 35982 15750 36034 15802
rect 36046 15750 36098 15802
rect 36110 15750 36162 15802
rect 66574 15750 66626 15802
rect 66638 15750 66690 15802
rect 66702 15750 66754 15802
rect 66766 15750 66818 15802
rect 66830 15750 66882 15802
rect 5794 15206 5846 15258
rect 5858 15206 5910 15258
rect 5922 15206 5974 15258
rect 5986 15206 6038 15258
rect 6050 15206 6102 15258
rect 36514 15206 36566 15258
rect 36578 15206 36630 15258
rect 36642 15206 36694 15258
rect 36706 15206 36758 15258
rect 36770 15206 36822 15258
rect 67234 15206 67286 15258
rect 67298 15206 67350 15258
rect 67362 15206 67414 15258
rect 67426 15206 67478 15258
rect 67490 15206 67542 15258
rect 5134 14662 5186 14714
rect 5198 14662 5250 14714
rect 5262 14662 5314 14714
rect 5326 14662 5378 14714
rect 5390 14662 5442 14714
rect 35854 14662 35906 14714
rect 35918 14662 35970 14714
rect 35982 14662 36034 14714
rect 36046 14662 36098 14714
rect 36110 14662 36162 14714
rect 66574 14662 66626 14714
rect 66638 14662 66690 14714
rect 66702 14662 66754 14714
rect 66766 14662 66818 14714
rect 66830 14662 66882 14714
rect 5794 14118 5846 14170
rect 5858 14118 5910 14170
rect 5922 14118 5974 14170
rect 5986 14118 6038 14170
rect 6050 14118 6102 14170
rect 36514 14118 36566 14170
rect 36578 14118 36630 14170
rect 36642 14118 36694 14170
rect 36706 14118 36758 14170
rect 36770 14118 36822 14170
rect 67234 14118 67286 14170
rect 67298 14118 67350 14170
rect 67362 14118 67414 14170
rect 67426 14118 67478 14170
rect 67490 14118 67542 14170
rect 5134 13574 5186 13626
rect 5198 13574 5250 13626
rect 5262 13574 5314 13626
rect 5326 13574 5378 13626
rect 5390 13574 5442 13626
rect 35854 13574 35906 13626
rect 35918 13574 35970 13626
rect 35982 13574 36034 13626
rect 36046 13574 36098 13626
rect 36110 13574 36162 13626
rect 66574 13574 66626 13626
rect 66638 13574 66690 13626
rect 66702 13574 66754 13626
rect 66766 13574 66818 13626
rect 66830 13574 66882 13626
rect 5794 13030 5846 13082
rect 5858 13030 5910 13082
rect 5922 13030 5974 13082
rect 5986 13030 6038 13082
rect 6050 13030 6102 13082
rect 36514 13030 36566 13082
rect 36578 13030 36630 13082
rect 36642 13030 36694 13082
rect 36706 13030 36758 13082
rect 36770 13030 36822 13082
rect 67234 13030 67286 13082
rect 67298 13030 67350 13082
rect 67362 13030 67414 13082
rect 67426 13030 67478 13082
rect 67490 13030 67542 13082
rect 5134 12486 5186 12538
rect 5198 12486 5250 12538
rect 5262 12486 5314 12538
rect 5326 12486 5378 12538
rect 5390 12486 5442 12538
rect 35854 12486 35906 12538
rect 35918 12486 35970 12538
rect 35982 12486 36034 12538
rect 36046 12486 36098 12538
rect 36110 12486 36162 12538
rect 66574 12486 66626 12538
rect 66638 12486 66690 12538
rect 66702 12486 66754 12538
rect 66766 12486 66818 12538
rect 66830 12486 66882 12538
rect 5794 11942 5846 11994
rect 5858 11942 5910 11994
rect 5922 11942 5974 11994
rect 5986 11942 6038 11994
rect 6050 11942 6102 11994
rect 36514 11942 36566 11994
rect 36578 11942 36630 11994
rect 36642 11942 36694 11994
rect 36706 11942 36758 11994
rect 36770 11942 36822 11994
rect 67234 11942 67286 11994
rect 67298 11942 67350 11994
rect 67362 11942 67414 11994
rect 67426 11942 67478 11994
rect 67490 11942 67542 11994
rect 5134 11398 5186 11450
rect 5198 11398 5250 11450
rect 5262 11398 5314 11450
rect 5326 11398 5378 11450
rect 5390 11398 5442 11450
rect 35854 11398 35906 11450
rect 35918 11398 35970 11450
rect 35982 11398 36034 11450
rect 36046 11398 36098 11450
rect 36110 11398 36162 11450
rect 66574 11398 66626 11450
rect 66638 11398 66690 11450
rect 66702 11398 66754 11450
rect 66766 11398 66818 11450
rect 66830 11398 66882 11450
rect 5794 10854 5846 10906
rect 5858 10854 5910 10906
rect 5922 10854 5974 10906
rect 5986 10854 6038 10906
rect 6050 10854 6102 10906
rect 36514 10854 36566 10906
rect 36578 10854 36630 10906
rect 36642 10854 36694 10906
rect 36706 10854 36758 10906
rect 36770 10854 36822 10906
rect 67234 10854 67286 10906
rect 67298 10854 67350 10906
rect 67362 10854 67414 10906
rect 67426 10854 67478 10906
rect 67490 10854 67542 10906
rect 5134 10310 5186 10362
rect 5198 10310 5250 10362
rect 5262 10310 5314 10362
rect 5326 10310 5378 10362
rect 5390 10310 5442 10362
rect 35854 10310 35906 10362
rect 35918 10310 35970 10362
rect 35982 10310 36034 10362
rect 36046 10310 36098 10362
rect 36110 10310 36162 10362
rect 66574 10310 66626 10362
rect 66638 10310 66690 10362
rect 66702 10310 66754 10362
rect 66766 10310 66818 10362
rect 66830 10310 66882 10362
rect 5794 9766 5846 9818
rect 5858 9766 5910 9818
rect 5922 9766 5974 9818
rect 5986 9766 6038 9818
rect 6050 9766 6102 9818
rect 36514 9766 36566 9818
rect 36578 9766 36630 9818
rect 36642 9766 36694 9818
rect 36706 9766 36758 9818
rect 36770 9766 36822 9818
rect 67234 9766 67286 9818
rect 67298 9766 67350 9818
rect 67362 9766 67414 9818
rect 67426 9766 67478 9818
rect 67490 9766 67542 9818
rect 5134 9222 5186 9274
rect 5198 9222 5250 9274
rect 5262 9222 5314 9274
rect 5326 9222 5378 9274
rect 5390 9222 5442 9274
rect 35854 9222 35906 9274
rect 35918 9222 35970 9274
rect 35982 9222 36034 9274
rect 36046 9222 36098 9274
rect 36110 9222 36162 9274
rect 66574 9222 66626 9274
rect 66638 9222 66690 9274
rect 66702 9222 66754 9274
rect 66766 9222 66818 9274
rect 66830 9222 66882 9274
rect 5794 8678 5846 8730
rect 5858 8678 5910 8730
rect 5922 8678 5974 8730
rect 5986 8678 6038 8730
rect 6050 8678 6102 8730
rect 36514 8678 36566 8730
rect 36578 8678 36630 8730
rect 36642 8678 36694 8730
rect 36706 8678 36758 8730
rect 36770 8678 36822 8730
rect 67234 8678 67286 8730
rect 67298 8678 67350 8730
rect 67362 8678 67414 8730
rect 67426 8678 67478 8730
rect 67490 8678 67542 8730
rect 5134 8134 5186 8186
rect 5198 8134 5250 8186
rect 5262 8134 5314 8186
rect 5326 8134 5378 8186
rect 5390 8134 5442 8186
rect 35854 8134 35906 8186
rect 35918 8134 35970 8186
rect 35982 8134 36034 8186
rect 36046 8134 36098 8186
rect 36110 8134 36162 8186
rect 66574 8134 66626 8186
rect 66638 8134 66690 8186
rect 66702 8134 66754 8186
rect 66766 8134 66818 8186
rect 66830 8134 66882 8186
rect 5794 7590 5846 7642
rect 5858 7590 5910 7642
rect 5922 7590 5974 7642
rect 5986 7590 6038 7642
rect 6050 7590 6102 7642
rect 36514 7590 36566 7642
rect 36578 7590 36630 7642
rect 36642 7590 36694 7642
rect 36706 7590 36758 7642
rect 36770 7590 36822 7642
rect 67234 7590 67286 7642
rect 67298 7590 67350 7642
rect 67362 7590 67414 7642
rect 67426 7590 67478 7642
rect 67490 7590 67542 7642
rect 5134 7046 5186 7098
rect 5198 7046 5250 7098
rect 5262 7046 5314 7098
rect 5326 7046 5378 7098
rect 5390 7046 5442 7098
rect 35854 7046 35906 7098
rect 35918 7046 35970 7098
rect 35982 7046 36034 7098
rect 36046 7046 36098 7098
rect 36110 7046 36162 7098
rect 66574 7046 66626 7098
rect 66638 7046 66690 7098
rect 66702 7046 66754 7098
rect 66766 7046 66818 7098
rect 66830 7046 66882 7098
rect 5794 6502 5846 6554
rect 5858 6502 5910 6554
rect 5922 6502 5974 6554
rect 5986 6502 6038 6554
rect 6050 6502 6102 6554
rect 36514 6502 36566 6554
rect 36578 6502 36630 6554
rect 36642 6502 36694 6554
rect 36706 6502 36758 6554
rect 36770 6502 36822 6554
rect 67234 6502 67286 6554
rect 67298 6502 67350 6554
rect 67362 6502 67414 6554
rect 67426 6502 67478 6554
rect 67490 6502 67542 6554
rect 5134 5958 5186 6010
rect 5198 5958 5250 6010
rect 5262 5958 5314 6010
rect 5326 5958 5378 6010
rect 5390 5958 5442 6010
rect 35854 5958 35906 6010
rect 35918 5958 35970 6010
rect 35982 5958 36034 6010
rect 36046 5958 36098 6010
rect 36110 5958 36162 6010
rect 66574 5958 66626 6010
rect 66638 5958 66690 6010
rect 66702 5958 66754 6010
rect 66766 5958 66818 6010
rect 66830 5958 66882 6010
rect 5794 5414 5846 5466
rect 5858 5414 5910 5466
rect 5922 5414 5974 5466
rect 5986 5414 6038 5466
rect 6050 5414 6102 5466
rect 36514 5414 36566 5466
rect 36578 5414 36630 5466
rect 36642 5414 36694 5466
rect 36706 5414 36758 5466
rect 36770 5414 36822 5466
rect 67234 5414 67286 5466
rect 67298 5414 67350 5466
rect 67362 5414 67414 5466
rect 67426 5414 67478 5466
rect 67490 5414 67542 5466
rect 5134 4870 5186 4922
rect 5198 4870 5250 4922
rect 5262 4870 5314 4922
rect 5326 4870 5378 4922
rect 5390 4870 5442 4922
rect 35854 4870 35906 4922
rect 35918 4870 35970 4922
rect 35982 4870 36034 4922
rect 36046 4870 36098 4922
rect 36110 4870 36162 4922
rect 66574 4870 66626 4922
rect 66638 4870 66690 4922
rect 66702 4870 66754 4922
rect 66766 4870 66818 4922
rect 66830 4870 66882 4922
rect 5794 4326 5846 4378
rect 5858 4326 5910 4378
rect 5922 4326 5974 4378
rect 5986 4326 6038 4378
rect 6050 4326 6102 4378
rect 36514 4326 36566 4378
rect 36578 4326 36630 4378
rect 36642 4326 36694 4378
rect 36706 4326 36758 4378
rect 36770 4326 36822 4378
rect 67234 4326 67286 4378
rect 67298 4326 67350 4378
rect 67362 4326 67414 4378
rect 67426 4326 67478 4378
rect 67490 4326 67542 4378
rect 5134 3782 5186 3834
rect 5198 3782 5250 3834
rect 5262 3782 5314 3834
rect 5326 3782 5378 3834
rect 5390 3782 5442 3834
rect 35854 3782 35906 3834
rect 35918 3782 35970 3834
rect 35982 3782 36034 3834
rect 36046 3782 36098 3834
rect 36110 3782 36162 3834
rect 66574 3782 66626 3834
rect 66638 3782 66690 3834
rect 66702 3782 66754 3834
rect 66766 3782 66818 3834
rect 66830 3782 66882 3834
rect 5794 3238 5846 3290
rect 5858 3238 5910 3290
rect 5922 3238 5974 3290
rect 5986 3238 6038 3290
rect 6050 3238 6102 3290
rect 36514 3238 36566 3290
rect 36578 3238 36630 3290
rect 36642 3238 36694 3290
rect 36706 3238 36758 3290
rect 36770 3238 36822 3290
rect 67234 3238 67286 3290
rect 67298 3238 67350 3290
rect 67362 3238 67414 3290
rect 67426 3238 67478 3290
rect 67490 3238 67542 3290
rect 5134 2694 5186 2746
rect 5198 2694 5250 2746
rect 5262 2694 5314 2746
rect 5326 2694 5378 2746
rect 5390 2694 5442 2746
rect 35854 2694 35906 2746
rect 35918 2694 35970 2746
rect 35982 2694 36034 2746
rect 36046 2694 36098 2746
rect 36110 2694 36162 2746
rect 66574 2694 66626 2746
rect 66638 2694 66690 2746
rect 66702 2694 66754 2746
rect 66766 2694 66818 2746
rect 66830 2694 66882 2746
rect 22560 2388 22612 2440
rect 23204 2388 23256 2440
rect 33508 2388 33560 2440
rect 41880 2388 41932 2440
rect 42524 2388 42576 2440
rect 44456 2388 44508 2440
rect 52184 2388 52236 2440
rect 57980 2388 58032 2440
rect 59268 2388 59320 2440
rect 5794 2150 5846 2202
rect 5858 2150 5910 2202
rect 5922 2150 5974 2202
rect 5986 2150 6038 2202
rect 6050 2150 6102 2202
rect 36514 2150 36566 2202
rect 36578 2150 36630 2202
rect 36642 2150 36694 2202
rect 36706 2150 36758 2202
rect 36770 2150 36822 2202
rect 67234 2150 67286 2202
rect 67298 2150 67350 2202
rect 67362 2150 67414 2202
rect 67426 2150 67478 2202
rect 67490 2150 67542 2202
<< metal2 >>
rect 23846 79200 23902 80000
rect 32862 79200 32918 80000
rect 39946 79200 40002 80000
rect 41878 79200 41934 80000
rect 49606 79200 49662 80000
rect 54114 79200 54170 80000
rect 58622 79200 58678 80000
rect 5134 77820 5442 77829
rect 5134 77818 5140 77820
rect 5196 77818 5220 77820
rect 5276 77818 5300 77820
rect 5356 77818 5380 77820
rect 5436 77818 5442 77820
rect 5196 77766 5198 77818
rect 5378 77766 5380 77818
rect 5134 77764 5140 77766
rect 5196 77764 5220 77766
rect 5276 77764 5300 77766
rect 5356 77764 5380 77766
rect 5436 77764 5442 77766
rect 5134 77755 5442 77764
rect 23860 77722 23888 79200
rect 32876 77722 32904 79200
rect 35854 77820 36162 77829
rect 35854 77818 35860 77820
rect 35916 77818 35940 77820
rect 35996 77818 36020 77820
rect 36076 77818 36100 77820
rect 36156 77818 36162 77820
rect 35916 77766 35918 77818
rect 36098 77766 36100 77818
rect 35854 77764 35860 77766
rect 35916 77764 35940 77766
rect 35996 77764 36020 77766
rect 36076 77764 36100 77766
rect 36156 77764 36162 77766
rect 35854 77755 36162 77764
rect 39960 77722 39988 79200
rect 41892 77722 41920 79200
rect 49620 77722 49648 79200
rect 54128 77722 54156 79200
rect 58636 77722 58664 79200
rect 66574 77820 66882 77829
rect 66574 77818 66580 77820
rect 66636 77818 66660 77820
rect 66716 77818 66740 77820
rect 66796 77818 66820 77820
rect 66876 77818 66882 77820
rect 66636 77766 66638 77818
rect 66818 77766 66820 77818
rect 66574 77764 66580 77766
rect 66636 77764 66660 77766
rect 66716 77764 66740 77766
rect 66796 77764 66820 77766
rect 66876 77764 66882 77766
rect 66574 77755 66882 77764
rect 23848 77716 23900 77722
rect 23848 77658 23900 77664
rect 32864 77716 32916 77722
rect 32864 77658 32916 77664
rect 39948 77716 40000 77722
rect 39948 77658 40000 77664
rect 41880 77716 41932 77722
rect 41880 77658 41932 77664
rect 49608 77716 49660 77722
rect 49608 77658 49660 77664
rect 54116 77716 54168 77722
rect 54116 77658 54168 77664
rect 58624 77716 58676 77722
rect 58624 77658 58676 77664
rect 5794 77276 6102 77285
rect 5794 77274 5800 77276
rect 5856 77274 5880 77276
rect 5936 77274 5960 77276
rect 6016 77274 6040 77276
rect 6096 77274 6102 77276
rect 5856 77222 5858 77274
rect 6038 77222 6040 77274
rect 5794 77220 5800 77222
rect 5856 77220 5880 77222
rect 5936 77220 5960 77222
rect 6016 77220 6040 77222
rect 6096 77220 6102 77222
rect 5794 77211 6102 77220
rect 36514 77276 36822 77285
rect 36514 77274 36520 77276
rect 36576 77274 36600 77276
rect 36656 77274 36680 77276
rect 36736 77274 36760 77276
rect 36816 77274 36822 77276
rect 36576 77222 36578 77274
rect 36758 77222 36760 77274
rect 36514 77220 36520 77222
rect 36576 77220 36600 77222
rect 36656 77220 36680 77222
rect 36736 77220 36760 77222
rect 36816 77220 36822 77222
rect 36514 77211 36822 77220
rect 67234 77276 67542 77285
rect 67234 77274 67240 77276
rect 67296 77274 67320 77276
rect 67376 77274 67400 77276
rect 67456 77274 67480 77276
rect 67536 77274 67542 77276
rect 67296 77222 67298 77274
rect 67478 77222 67480 77274
rect 67234 77220 67240 77222
rect 67296 77220 67320 77222
rect 67376 77220 67400 77222
rect 67456 77220 67480 77222
rect 67536 77220 67542 77222
rect 67234 77211 67542 77220
rect 5134 76732 5442 76741
rect 5134 76730 5140 76732
rect 5196 76730 5220 76732
rect 5276 76730 5300 76732
rect 5356 76730 5380 76732
rect 5436 76730 5442 76732
rect 5196 76678 5198 76730
rect 5378 76678 5380 76730
rect 5134 76676 5140 76678
rect 5196 76676 5220 76678
rect 5276 76676 5300 76678
rect 5356 76676 5380 76678
rect 5436 76676 5442 76678
rect 5134 76667 5442 76676
rect 35854 76732 36162 76741
rect 35854 76730 35860 76732
rect 35916 76730 35940 76732
rect 35996 76730 36020 76732
rect 36076 76730 36100 76732
rect 36156 76730 36162 76732
rect 35916 76678 35918 76730
rect 36098 76678 36100 76730
rect 35854 76676 35860 76678
rect 35916 76676 35940 76678
rect 35996 76676 36020 76678
rect 36076 76676 36100 76678
rect 36156 76676 36162 76678
rect 35854 76667 36162 76676
rect 66574 76732 66882 76741
rect 66574 76730 66580 76732
rect 66636 76730 66660 76732
rect 66716 76730 66740 76732
rect 66796 76730 66820 76732
rect 66876 76730 66882 76732
rect 66636 76678 66638 76730
rect 66818 76678 66820 76730
rect 66574 76676 66580 76678
rect 66636 76676 66660 76678
rect 66716 76676 66740 76678
rect 66796 76676 66820 76678
rect 66876 76676 66882 76678
rect 66574 76667 66882 76676
rect 5794 76188 6102 76197
rect 5794 76186 5800 76188
rect 5856 76186 5880 76188
rect 5936 76186 5960 76188
rect 6016 76186 6040 76188
rect 6096 76186 6102 76188
rect 5856 76134 5858 76186
rect 6038 76134 6040 76186
rect 5794 76132 5800 76134
rect 5856 76132 5880 76134
rect 5936 76132 5960 76134
rect 6016 76132 6040 76134
rect 6096 76132 6102 76134
rect 5794 76123 6102 76132
rect 36514 76188 36822 76197
rect 36514 76186 36520 76188
rect 36576 76186 36600 76188
rect 36656 76186 36680 76188
rect 36736 76186 36760 76188
rect 36816 76186 36822 76188
rect 36576 76134 36578 76186
rect 36758 76134 36760 76186
rect 36514 76132 36520 76134
rect 36576 76132 36600 76134
rect 36656 76132 36680 76134
rect 36736 76132 36760 76134
rect 36816 76132 36822 76134
rect 36514 76123 36822 76132
rect 67234 76188 67542 76197
rect 67234 76186 67240 76188
rect 67296 76186 67320 76188
rect 67376 76186 67400 76188
rect 67456 76186 67480 76188
rect 67536 76186 67542 76188
rect 67296 76134 67298 76186
rect 67478 76134 67480 76186
rect 67234 76132 67240 76134
rect 67296 76132 67320 76134
rect 67376 76132 67400 76134
rect 67456 76132 67480 76134
rect 67536 76132 67542 76134
rect 67234 76123 67542 76132
rect 5134 75644 5442 75653
rect 5134 75642 5140 75644
rect 5196 75642 5220 75644
rect 5276 75642 5300 75644
rect 5356 75642 5380 75644
rect 5436 75642 5442 75644
rect 5196 75590 5198 75642
rect 5378 75590 5380 75642
rect 5134 75588 5140 75590
rect 5196 75588 5220 75590
rect 5276 75588 5300 75590
rect 5356 75588 5380 75590
rect 5436 75588 5442 75590
rect 5134 75579 5442 75588
rect 35854 75644 36162 75653
rect 35854 75642 35860 75644
rect 35916 75642 35940 75644
rect 35996 75642 36020 75644
rect 36076 75642 36100 75644
rect 36156 75642 36162 75644
rect 35916 75590 35918 75642
rect 36098 75590 36100 75642
rect 35854 75588 35860 75590
rect 35916 75588 35940 75590
rect 35996 75588 36020 75590
rect 36076 75588 36100 75590
rect 36156 75588 36162 75590
rect 35854 75579 36162 75588
rect 66574 75644 66882 75653
rect 66574 75642 66580 75644
rect 66636 75642 66660 75644
rect 66716 75642 66740 75644
rect 66796 75642 66820 75644
rect 66876 75642 66882 75644
rect 66636 75590 66638 75642
rect 66818 75590 66820 75642
rect 66574 75588 66580 75590
rect 66636 75588 66660 75590
rect 66716 75588 66740 75590
rect 66796 75588 66820 75590
rect 66876 75588 66882 75590
rect 66574 75579 66882 75588
rect 5794 75100 6102 75109
rect 5794 75098 5800 75100
rect 5856 75098 5880 75100
rect 5936 75098 5960 75100
rect 6016 75098 6040 75100
rect 6096 75098 6102 75100
rect 5856 75046 5858 75098
rect 6038 75046 6040 75098
rect 5794 75044 5800 75046
rect 5856 75044 5880 75046
rect 5936 75044 5960 75046
rect 6016 75044 6040 75046
rect 6096 75044 6102 75046
rect 5794 75035 6102 75044
rect 36514 75100 36822 75109
rect 36514 75098 36520 75100
rect 36576 75098 36600 75100
rect 36656 75098 36680 75100
rect 36736 75098 36760 75100
rect 36816 75098 36822 75100
rect 36576 75046 36578 75098
rect 36758 75046 36760 75098
rect 36514 75044 36520 75046
rect 36576 75044 36600 75046
rect 36656 75044 36680 75046
rect 36736 75044 36760 75046
rect 36816 75044 36822 75046
rect 36514 75035 36822 75044
rect 67234 75100 67542 75109
rect 67234 75098 67240 75100
rect 67296 75098 67320 75100
rect 67376 75098 67400 75100
rect 67456 75098 67480 75100
rect 67536 75098 67542 75100
rect 67296 75046 67298 75098
rect 67478 75046 67480 75098
rect 67234 75044 67240 75046
rect 67296 75044 67320 75046
rect 67376 75044 67400 75046
rect 67456 75044 67480 75046
rect 67536 75044 67542 75046
rect 67234 75035 67542 75044
rect 5134 74556 5442 74565
rect 5134 74554 5140 74556
rect 5196 74554 5220 74556
rect 5276 74554 5300 74556
rect 5356 74554 5380 74556
rect 5436 74554 5442 74556
rect 5196 74502 5198 74554
rect 5378 74502 5380 74554
rect 5134 74500 5140 74502
rect 5196 74500 5220 74502
rect 5276 74500 5300 74502
rect 5356 74500 5380 74502
rect 5436 74500 5442 74502
rect 5134 74491 5442 74500
rect 35854 74556 36162 74565
rect 35854 74554 35860 74556
rect 35916 74554 35940 74556
rect 35996 74554 36020 74556
rect 36076 74554 36100 74556
rect 36156 74554 36162 74556
rect 35916 74502 35918 74554
rect 36098 74502 36100 74554
rect 35854 74500 35860 74502
rect 35916 74500 35940 74502
rect 35996 74500 36020 74502
rect 36076 74500 36100 74502
rect 36156 74500 36162 74502
rect 35854 74491 36162 74500
rect 66574 74556 66882 74565
rect 66574 74554 66580 74556
rect 66636 74554 66660 74556
rect 66716 74554 66740 74556
rect 66796 74554 66820 74556
rect 66876 74554 66882 74556
rect 66636 74502 66638 74554
rect 66818 74502 66820 74554
rect 66574 74500 66580 74502
rect 66636 74500 66660 74502
rect 66716 74500 66740 74502
rect 66796 74500 66820 74502
rect 66876 74500 66882 74502
rect 66574 74491 66882 74500
rect 5794 74012 6102 74021
rect 5794 74010 5800 74012
rect 5856 74010 5880 74012
rect 5936 74010 5960 74012
rect 6016 74010 6040 74012
rect 6096 74010 6102 74012
rect 5856 73958 5858 74010
rect 6038 73958 6040 74010
rect 5794 73956 5800 73958
rect 5856 73956 5880 73958
rect 5936 73956 5960 73958
rect 6016 73956 6040 73958
rect 6096 73956 6102 73958
rect 5794 73947 6102 73956
rect 36514 74012 36822 74021
rect 36514 74010 36520 74012
rect 36576 74010 36600 74012
rect 36656 74010 36680 74012
rect 36736 74010 36760 74012
rect 36816 74010 36822 74012
rect 36576 73958 36578 74010
rect 36758 73958 36760 74010
rect 36514 73956 36520 73958
rect 36576 73956 36600 73958
rect 36656 73956 36680 73958
rect 36736 73956 36760 73958
rect 36816 73956 36822 73958
rect 36514 73947 36822 73956
rect 67234 74012 67542 74021
rect 67234 74010 67240 74012
rect 67296 74010 67320 74012
rect 67376 74010 67400 74012
rect 67456 74010 67480 74012
rect 67536 74010 67542 74012
rect 67296 73958 67298 74010
rect 67478 73958 67480 74010
rect 67234 73956 67240 73958
rect 67296 73956 67320 73958
rect 67376 73956 67400 73958
rect 67456 73956 67480 73958
rect 67536 73956 67542 73958
rect 67234 73947 67542 73956
rect 5134 73468 5442 73477
rect 5134 73466 5140 73468
rect 5196 73466 5220 73468
rect 5276 73466 5300 73468
rect 5356 73466 5380 73468
rect 5436 73466 5442 73468
rect 5196 73414 5198 73466
rect 5378 73414 5380 73466
rect 5134 73412 5140 73414
rect 5196 73412 5220 73414
rect 5276 73412 5300 73414
rect 5356 73412 5380 73414
rect 5436 73412 5442 73414
rect 5134 73403 5442 73412
rect 35854 73468 36162 73477
rect 35854 73466 35860 73468
rect 35916 73466 35940 73468
rect 35996 73466 36020 73468
rect 36076 73466 36100 73468
rect 36156 73466 36162 73468
rect 35916 73414 35918 73466
rect 36098 73414 36100 73466
rect 35854 73412 35860 73414
rect 35916 73412 35940 73414
rect 35996 73412 36020 73414
rect 36076 73412 36100 73414
rect 36156 73412 36162 73414
rect 35854 73403 36162 73412
rect 66574 73468 66882 73477
rect 66574 73466 66580 73468
rect 66636 73466 66660 73468
rect 66716 73466 66740 73468
rect 66796 73466 66820 73468
rect 66876 73466 66882 73468
rect 66636 73414 66638 73466
rect 66818 73414 66820 73466
rect 66574 73412 66580 73414
rect 66636 73412 66660 73414
rect 66716 73412 66740 73414
rect 66796 73412 66820 73414
rect 66876 73412 66882 73414
rect 66574 73403 66882 73412
rect 5794 72924 6102 72933
rect 5794 72922 5800 72924
rect 5856 72922 5880 72924
rect 5936 72922 5960 72924
rect 6016 72922 6040 72924
rect 6096 72922 6102 72924
rect 5856 72870 5858 72922
rect 6038 72870 6040 72922
rect 5794 72868 5800 72870
rect 5856 72868 5880 72870
rect 5936 72868 5960 72870
rect 6016 72868 6040 72870
rect 6096 72868 6102 72870
rect 5794 72859 6102 72868
rect 36514 72924 36822 72933
rect 36514 72922 36520 72924
rect 36576 72922 36600 72924
rect 36656 72922 36680 72924
rect 36736 72922 36760 72924
rect 36816 72922 36822 72924
rect 36576 72870 36578 72922
rect 36758 72870 36760 72922
rect 36514 72868 36520 72870
rect 36576 72868 36600 72870
rect 36656 72868 36680 72870
rect 36736 72868 36760 72870
rect 36816 72868 36822 72870
rect 36514 72859 36822 72868
rect 67234 72924 67542 72933
rect 67234 72922 67240 72924
rect 67296 72922 67320 72924
rect 67376 72922 67400 72924
rect 67456 72922 67480 72924
rect 67536 72922 67542 72924
rect 67296 72870 67298 72922
rect 67478 72870 67480 72922
rect 67234 72868 67240 72870
rect 67296 72868 67320 72870
rect 67376 72868 67400 72870
rect 67456 72868 67480 72870
rect 67536 72868 67542 72870
rect 67234 72859 67542 72868
rect 5134 72380 5442 72389
rect 5134 72378 5140 72380
rect 5196 72378 5220 72380
rect 5276 72378 5300 72380
rect 5356 72378 5380 72380
rect 5436 72378 5442 72380
rect 5196 72326 5198 72378
rect 5378 72326 5380 72378
rect 5134 72324 5140 72326
rect 5196 72324 5220 72326
rect 5276 72324 5300 72326
rect 5356 72324 5380 72326
rect 5436 72324 5442 72326
rect 5134 72315 5442 72324
rect 35854 72380 36162 72389
rect 35854 72378 35860 72380
rect 35916 72378 35940 72380
rect 35996 72378 36020 72380
rect 36076 72378 36100 72380
rect 36156 72378 36162 72380
rect 35916 72326 35918 72378
rect 36098 72326 36100 72378
rect 35854 72324 35860 72326
rect 35916 72324 35940 72326
rect 35996 72324 36020 72326
rect 36076 72324 36100 72326
rect 36156 72324 36162 72326
rect 35854 72315 36162 72324
rect 66574 72380 66882 72389
rect 66574 72378 66580 72380
rect 66636 72378 66660 72380
rect 66716 72378 66740 72380
rect 66796 72378 66820 72380
rect 66876 72378 66882 72380
rect 66636 72326 66638 72378
rect 66818 72326 66820 72378
rect 66574 72324 66580 72326
rect 66636 72324 66660 72326
rect 66716 72324 66740 72326
rect 66796 72324 66820 72326
rect 66876 72324 66882 72326
rect 66574 72315 66882 72324
rect 5794 71836 6102 71845
rect 5794 71834 5800 71836
rect 5856 71834 5880 71836
rect 5936 71834 5960 71836
rect 6016 71834 6040 71836
rect 6096 71834 6102 71836
rect 5856 71782 5858 71834
rect 6038 71782 6040 71834
rect 5794 71780 5800 71782
rect 5856 71780 5880 71782
rect 5936 71780 5960 71782
rect 6016 71780 6040 71782
rect 6096 71780 6102 71782
rect 5794 71771 6102 71780
rect 36514 71836 36822 71845
rect 36514 71834 36520 71836
rect 36576 71834 36600 71836
rect 36656 71834 36680 71836
rect 36736 71834 36760 71836
rect 36816 71834 36822 71836
rect 36576 71782 36578 71834
rect 36758 71782 36760 71834
rect 36514 71780 36520 71782
rect 36576 71780 36600 71782
rect 36656 71780 36680 71782
rect 36736 71780 36760 71782
rect 36816 71780 36822 71782
rect 36514 71771 36822 71780
rect 67234 71836 67542 71845
rect 67234 71834 67240 71836
rect 67296 71834 67320 71836
rect 67376 71834 67400 71836
rect 67456 71834 67480 71836
rect 67536 71834 67542 71836
rect 67296 71782 67298 71834
rect 67478 71782 67480 71834
rect 67234 71780 67240 71782
rect 67296 71780 67320 71782
rect 67376 71780 67400 71782
rect 67456 71780 67480 71782
rect 67536 71780 67542 71782
rect 67234 71771 67542 71780
rect 5134 71292 5442 71301
rect 5134 71290 5140 71292
rect 5196 71290 5220 71292
rect 5276 71290 5300 71292
rect 5356 71290 5380 71292
rect 5436 71290 5442 71292
rect 5196 71238 5198 71290
rect 5378 71238 5380 71290
rect 5134 71236 5140 71238
rect 5196 71236 5220 71238
rect 5276 71236 5300 71238
rect 5356 71236 5380 71238
rect 5436 71236 5442 71238
rect 5134 71227 5442 71236
rect 35854 71292 36162 71301
rect 35854 71290 35860 71292
rect 35916 71290 35940 71292
rect 35996 71290 36020 71292
rect 36076 71290 36100 71292
rect 36156 71290 36162 71292
rect 35916 71238 35918 71290
rect 36098 71238 36100 71290
rect 35854 71236 35860 71238
rect 35916 71236 35940 71238
rect 35996 71236 36020 71238
rect 36076 71236 36100 71238
rect 36156 71236 36162 71238
rect 35854 71227 36162 71236
rect 66574 71292 66882 71301
rect 66574 71290 66580 71292
rect 66636 71290 66660 71292
rect 66716 71290 66740 71292
rect 66796 71290 66820 71292
rect 66876 71290 66882 71292
rect 66636 71238 66638 71290
rect 66818 71238 66820 71290
rect 66574 71236 66580 71238
rect 66636 71236 66660 71238
rect 66716 71236 66740 71238
rect 66796 71236 66820 71238
rect 66876 71236 66882 71238
rect 66574 71227 66882 71236
rect 5794 70748 6102 70757
rect 5794 70746 5800 70748
rect 5856 70746 5880 70748
rect 5936 70746 5960 70748
rect 6016 70746 6040 70748
rect 6096 70746 6102 70748
rect 5856 70694 5858 70746
rect 6038 70694 6040 70746
rect 5794 70692 5800 70694
rect 5856 70692 5880 70694
rect 5936 70692 5960 70694
rect 6016 70692 6040 70694
rect 6096 70692 6102 70694
rect 5794 70683 6102 70692
rect 36514 70748 36822 70757
rect 36514 70746 36520 70748
rect 36576 70746 36600 70748
rect 36656 70746 36680 70748
rect 36736 70746 36760 70748
rect 36816 70746 36822 70748
rect 36576 70694 36578 70746
rect 36758 70694 36760 70746
rect 36514 70692 36520 70694
rect 36576 70692 36600 70694
rect 36656 70692 36680 70694
rect 36736 70692 36760 70694
rect 36816 70692 36822 70694
rect 36514 70683 36822 70692
rect 67234 70748 67542 70757
rect 67234 70746 67240 70748
rect 67296 70746 67320 70748
rect 67376 70746 67400 70748
rect 67456 70746 67480 70748
rect 67536 70746 67542 70748
rect 67296 70694 67298 70746
rect 67478 70694 67480 70746
rect 67234 70692 67240 70694
rect 67296 70692 67320 70694
rect 67376 70692 67400 70694
rect 67456 70692 67480 70694
rect 67536 70692 67542 70694
rect 67234 70683 67542 70692
rect 5134 70204 5442 70213
rect 5134 70202 5140 70204
rect 5196 70202 5220 70204
rect 5276 70202 5300 70204
rect 5356 70202 5380 70204
rect 5436 70202 5442 70204
rect 5196 70150 5198 70202
rect 5378 70150 5380 70202
rect 5134 70148 5140 70150
rect 5196 70148 5220 70150
rect 5276 70148 5300 70150
rect 5356 70148 5380 70150
rect 5436 70148 5442 70150
rect 5134 70139 5442 70148
rect 35854 70204 36162 70213
rect 35854 70202 35860 70204
rect 35916 70202 35940 70204
rect 35996 70202 36020 70204
rect 36076 70202 36100 70204
rect 36156 70202 36162 70204
rect 35916 70150 35918 70202
rect 36098 70150 36100 70202
rect 35854 70148 35860 70150
rect 35916 70148 35940 70150
rect 35996 70148 36020 70150
rect 36076 70148 36100 70150
rect 36156 70148 36162 70150
rect 35854 70139 36162 70148
rect 66574 70204 66882 70213
rect 66574 70202 66580 70204
rect 66636 70202 66660 70204
rect 66716 70202 66740 70204
rect 66796 70202 66820 70204
rect 66876 70202 66882 70204
rect 66636 70150 66638 70202
rect 66818 70150 66820 70202
rect 66574 70148 66580 70150
rect 66636 70148 66660 70150
rect 66716 70148 66740 70150
rect 66796 70148 66820 70150
rect 66876 70148 66882 70150
rect 66574 70139 66882 70148
rect 5794 69660 6102 69669
rect 5794 69658 5800 69660
rect 5856 69658 5880 69660
rect 5936 69658 5960 69660
rect 6016 69658 6040 69660
rect 6096 69658 6102 69660
rect 5856 69606 5858 69658
rect 6038 69606 6040 69658
rect 5794 69604 5800 69606
rect 5856 69604 5880 69606
rect 5936 69604 5960 69606
rect 6016 69604 6040 69606
rect 6096 69604 6102 69606
rect 5794 69595 6102 69604
rect 36514 69660 36822 69669
rect 36514 69658 36520 69660
rect 36576 69658 36600 69660
rect 36656 69658 36680 69660
rect 36736 69658 36760 69660
rect 36816 69658 36822 69660
rect 36576 69606 36578 69658
rect 36758 69606 36760 69658
rect 36514 69604 36520 69606
rect 36576 69604 36600 69606
rect 36656 69604 36680 69606
rect 36736 69604 36760 69606
rect 36816 69604 36822 69606
rect 36514 69595 36822 69604
rect 67234 69660 67542 69669
rect 67234 69658 67240 69660
rect 67296 69658 67320 69660
rect 67376 69658 67400 69660
rect 67456 69658 67480 69660
rect 67536 69658 67542 69660
rect 67296 69606 67298 69658
rect 67478 69606 67480 69658
rect 67234 69604 67240 69606
rect 67296 69604 67320 69606
rect 67376 69604 67400 69606
rect 67456 69604 67480 69606
rect 67536 69604 67542 69606
rect 67234 69595 67542 69604
rect 5134 69116 5442 69125
rect 5134 69114 5140 69116
rect 5196 69114 5220 69116
rect 5276 69114 5300 69116
rect 5356 69114 5380 69116
rect 5436 69114 5442 69116
rect 5196 69062 5198 69114
rect 5378 69062 5380 69114
rect 5134 69060 5140 69062
rect 5196 69060 5220 69062
rect 5276 69060 5300 69062
rect 5356 69060 5380 69062
rect 5436 69060 5442 69062
rect 5134 69051 5442 69060
rect 35854 69116 36162 69125
rect 35854 69114 35860 69116
rect 35916 69114 35940 69116
rect 35996 69114 36020 69116
rect 36076 69114 36100 69116
rect 36156 69114 36162 69116
rect 35916 69062 35918 69114
rect 36098 69062 36100 69114
rect 35854 69060 35860 69062
rect 35916 69060 35940 69062
rect 35996 69060 36020 69062
rect 36076 69060 36100 69062
rect 36156 69060 36162 69062
rect 35854 69051 36162 69060
rect 66574 69116 66882 69125
rect 66574 69114 66580 69116
rect 66636 69114 66660 69116
rect 66716 69114 66740 69116
rect 66796 69114 66820 69116
rect 66876 69114 66882 69116
rect 66636 69062 66638 69114
rect 66818 69062 66820 69114
rect 66574 69060 66580 69062
rect 66636 69060 66660 69062
rect 66716 69060 66740 69062
rect 66796 69060 66820 69062
rect 66876 69060 66882 69062
rect 66574 69051 66882 69060
rect 5794 68572 6102 68581
rect 5794 68570 5800 68572
rect 5856 68570 5880 68572
rect 5936 68570 5960 68572
rect 6016 68570 6040 68572
rect 6096 68570 6102 68572
rect 5856 68518 5858 68570
rect 6038 68518 6040 68570
rect 5794 68516 5800 68518
rect 5856 68516 5880 68518
rect 5936 68516 5960 68518
rect 6016 68516 6040 68518
rect 6096 68516 6102 68518
rect 5794 68507 6102 68516
rect 36514 68572 36822 68581
rect 36514 68570 36520 68572
rect 36576 68570 36600 68572
rect 36656 68570 36680 68572
rect 36736 68570 36760 68572
rect 36816 68570 36822 68572
rect 36576 68518 36578 68570
rect 36758 68518 36760 68570
rect 36514 68516 36520 68518
rect 36576 68516 36600 68518
rect 36656 68516 36680 68518
rect 36736 68516 36760 68518
rect 36816 68516 36822 68518
rect 36514 68507 36822 68516
rect 67234 68572 67542 68581
rect 67234 68570 67240 68572
rect 67296 68570 67320 68572
rect 67376 68570 67400 68572
rect 67456 68570 67480 68572
rect 67536 68570 67542 68572
rect 67296 68518 67298 68570
rect 67478 68518 67480 68570
rect 67234 68516 67240 68518
rect 67296 68516 67320 68518
rect 67376 68516 67400 68518
rect 67456 68516 67480 68518
rect 67536 68516 67542 68518
rect 67234 68507 67542 68516
rect 5134 68028 5442 68037
rect 5134 68026 5140 68028
rect 5196 68026 5220 68028
rect 5276 68026 5300 68028
rect 5356 68026 5380 68028
rect 5436 68026 5442 68028
rect 5196 67974 5198 68026
rect 5378 67974 5380 68026
rect 5134 67972 5140 67974
rect 5196 67972 5220 67974
rect 5276 67972 5300 67974
rect 5356 67972 5380 67974
rect 5436 67972 5442 67974
rect 5134 67963 5442 67972
rect 35854 68028 36162 68037
rect 35854 68026 35860 68028
rect 35916 68026 35940 68028
rect 35996 68026 36020 68028
rect 36076 68026 36100 68028
rect 36156 68026 36162 68028
rect 35916 67974 35918 68026
rect 36098 67974 36100 68026
rect 35854 67972 35860 67974
rect 35916 67972 35940 67974
rect 35996 67972 36020 67974
rect 36076 67972 36100 67974
rect 36156 67972 36162 67974
rect 35854 67963 36162 67972
rect 66574 68028 66882 68037
rect 66574 68026 66580 68028
rect 66636 68026 66660 68028
rect 66716 68026 66740 68028
rect 66796 68026 66820 68028
rect 66876 68026 66882 68028
rect 66636 67974 66638 68026
rect 66818 67974 66820 68026
rect 66574 67972 66580 67974
rect 66636 67972 66660 67974
rect 66716 67972 66740 67974
rect 66796 67972 66820 67974
rect 66876 67972 66882 67974
rect 66574 67963 66882 67972
rect 5794 67484 6102 67493
rect 5794 67482 5800 67484
rect 5856 67482 5880 67484
rect 5936 67482 5960 67484
rect 6016 67482 6040 67484
rect 6096 67482 6102 67484
rect 5856 67430 5858 67482
rect 6038 67430 6040 67482
rect 5794 67428 5800 67430
rect 5856 67428 5880 67430
rect 5936 67428 5960 67430
rect 6016 67428 6040 67430
rect 6096 67428 6102 67430
rect 5794 67419 6102 67428
rect 36514 67484 36822 67493
rect 36514 67482 36520 67484
rect 36576 67482 36600 67484
rect 36656 67482 36680 67484
rect 36736 67482 36760 67484
rect 36816 67482 36822 67484
rect 36576 67430 36578 67482
rect 36758 67430 36760 67482
rect 36514 67428 36520 67430
rect 36576 67428 36600 67430
rect 36656 67428 36680 67430
rect 36736 67428 36760 67430
rect 36816 67428 36822 67430
rect 36514 67419 36822 67428
rect 67234 67484 67542 67493
rect 67234 67482 67240 67484
rect 67296 67482 67320 67484
rect 67376 67482 67400 67484
rect 67456 67482 67480 67484
rect 67536 67482 67542 67484
rect 67296 67430 67298 67482
rect 67478 67430 67480 67482
rect 67234 67428 67240 67430
rect 67296 67428 67320 67430
rect 67376 67428 67400 67430
rect 67456 67428 67480 67430
rect 67536 67428 67542 67430
rect 67234 67419 67542 67428
rect 5134 66940 5442 66949
rect 5134 66938 5140 66940
rect 5196 66938 5220 66940
rect 5276 66938 5300 66940
rect 5356 66938 5380 66940
rect 5436 66938 5442 66940
rect 5196 66886 5198 66938
rect 5378 66886 5380 66938
rect 5134 66884 5140 66886
rect 5196 66884 5220 66886
rect 5276 66884 5300 66886
rect 5356 66884 5380 66886
rect 5436 66884 5442 66886
rect 5134 66875 5442 66884
rect 35854 66940 36162 66949
rect 35854 66938 35860 66940
rect 35916 66938 35940 66940
rect 35996 66938 36020 66940
rect 36076 66938 36100 66940
rect 36156 66938 36162 66940
rect 35916 66886 35918 66938
rect 36098 66886 36100 66938
rect 35854 66884 35860 66886
rect 35916 66884 35940 66886
rect 35996 66884 36020 66886
rect 36076 66884 36100 66886
rect 36156 66884 36162 66886
rect 35854 66875 36162 66884
rect 66574 66940 66882 66949
rect 66574 66938 66580 66940
rect 66636 66938 66660 66940
rect 66716 66938 66740 66940
rect 66796 66938 66820 66940
rect 66876 66938 66882 66940
rect 66636 66886 66638 66938
rect 66818 66886 66820 66938
rect 66574 66884 66580 66886
rect 66636 66884 66660 66886
rect 66716 66884 66740 66886
rect 66796 66884 66820 66886
rect 66876 66884 66882 66886
rect 66574 66875 66882 66884
rect 5794 66396 6102 66405
rect 5794 66394 5800 66396
rect 5856 66394 5880 66396
rect 5936 66394 5960 66396
rect 6016 66394 6040 66396
rect 6096 66394 6102 66396
rect 5856 66342 5858 66394
rect 6038 66342 6040 66394
rect 5794 66340 5800 66342
rect 5856 66340 5880 66342
rect 5936 66340 5960 66342
rect 6016 66340 6040 66342
rect 6096 66340 6102 66342
rect 5794 66331 6102 66340
rect 36514 66396 36822 66405
rect 36514 66394 36520 66396
rect 36576 66394 36600 66396
rect 36656 66394 36680 66396
rect 36736 66394 36760 66396
rect 36816 66394 36822 66396
rect 36576 66342 36578 66394
rect 36758 66342 36760 66394
rect 36514 66340 36520 66342
rect 36576 66340 36600 66342
rect 36656 66340 36680 66342
rect 36736 66340 36760 66342
rect 36816 66340 36822 66342
rect 36514 66331 36822 66340
rect 67234 66396 67542 66405
rect 67234 66394 67240 66396
rect 67296 66394 67320 66396
rect 67376 66394 67400 66396
rect 67456 66394 67480 66396
rect 67536 66394 67542 66396
rect 67296 66342 67298 66394
rect 67478 66342 67480 66394
rect 67234 66340 67240 66342
rect 67296 66340 67320 66342
rect 67376 66340 67400 66342
rect 67456 66340 67480 66342
rect 67536 66340 67542 66342
rect 67234 66331 67542 66340
rect 5134 65852 5442 65861
rect 5134 65850 5140 65852
rect 5196 65850 5220 65852
rect 5276 65850 5300 65852
rect 5356 65850 5380 65852
rect 5436 65850 5442 65852
rect 5196 65798 5198 65850
rect 5378 65798 5380 65850
rect 5134 65796 5140 65798
rect 5196 65796 5220 65798
rect 5276 65796 5300 65798
rect 5356 65796 5380 65798
rect 5436 65796 5442 65798
rect 5134 65787 5442 65796
rect 35854 65852 36162 65861
rect 35854 65850 35860 65852
rect 35916 65850 35940 65852
rect 35996 65850 36020 65852
rect 36076 65850 36100 65852
rect 36156 65850 36162 65852
rect 35916 65798 35918 65850
rect 36098 65798 36100 65850
rect 35854 65796 35860 65798
rect 35916 65796 35940 65798
rect 35996 65796 36020 65798
rect 36076 65796 36100 65798
rect 36156 65796 36162 65798
rect 35854 65787 36162 65796
rect 66574 65852 66882 65861
rect 66574 65850 66580 65852
rect 66636 65850 66660 65852
rect 66716 65850 66740 65852
rect 66796 65850 66820 65852
rect 66876 65850 66882 65852
rect 66636 65798 66638 65850
rect 66818 65798 66820 65850
rect 66574 65796 66580 65798
rect 66636 65796 66660 65798
rect 66716 65796 66740 65798
rect 66796 65796 66820 65798
rect 66876 65796 66882 65798
rect 66574 65787 66882 65796
rect 5794 65308 6102 65317
rect 5794 65306 5800 65308
rect 5856 65306 5880 65308
rect 5936 65306 5960 65308
rect 6016 65306 6040 65308
rect 6096 65306 6102 65308
rect 5856 65254 5858 65306
rect 6038 65254 6040 65306
rect 5794 65252 5800 65254
rect 5856 65252 5880 65254
rect 5936 65252 5960 65254
rect 6016 65252 6040 65254
rect 6096 65252 6102 65254
rect 5794 65243 6102 65252
rect 36514 65308 36822 65317
rect 36514 65306 36520 65308
rect 36576 65306 36600 65308
rect 36656 65306 36680 65308
rect 36736 65306 36760 65308
rect 36816 65306 36822 65308
rect 36576 65254 36578 65306
rect 36758 65254 36760 65306
rect 36514 65252 36520 65254
rect 36576 65252 36600 65254
rect 36656 65252 36680 65254
rect 36736 65252 36760 65254
rect 36816 65252 36822 65254
rect 36514 65243 36822 65252
rect 67234 65308 67542 65317
rect 67234 65306 67240 65308
rect 67296 65306 67320 65308
rect 67376 65306 67400 65308
rect 67456 65306 67480 65308
rect 67536 65306 67542 65308
rect 67296 65254 67298 65306
rect 67478 65254 67480 65306
rect 67234 65252 67240 65254
rect 67296 65252 67320 65254
rect 67376 65252 67400 65254
rect 67456 65252 67480 65254
rect 67536 65252 67542 65254
rect 67234 65243 67542 65252
rect 5134 64764 5442 64773
rect 5134 64762 5140 64764
rect 5196 64762 5220 64764
rect 5276 64762 5300 64764
rect 5356 64762 5380 64764
rect 5436 64762 5442 64764
rect 5196 64710 5198 64762
rect 5378 64710 5380 64762
rect 5134 64708 5140 64710
rect 5196 64708 5220 64710
rect 5276 64708 5300 64710
rect 5356 64708 5380 64710
rect 5436 64708 5442 64710
rect 5134 64699 5442 64708
rect 35854 64764 36162 64773
rect 35854 64762 35860 64764
rect 35916 64762 35940 64764
rect 35996 64762 36020 64764
rect 36076 64762 36100 64764
rect 36156 64762 36162 64764
rect 35916 64710 35918 64762
rect 36098 64710 36100 64762
rect 35854 64708 35860 64710
rect 35916 64708 35940 64710
rect 35996 64708 36020 64710
rect 36076 64708 36100 64710
rect 36156 64708 36162 64710
rect 35854 64699 36162 64708
rect 66574 64764 66882 64773
rect 66574 64762 66580 64764
rect 66636 64762 66660 64764
rect 66716 64762 66740 64764
rect 66796 64762 66820 64764
rect 66876 64762 66882 64764
rect 66636 64710 66638 64762
rect 66818 64710 66820 64762
rect 66574 64708 66580 64710
rect 66636 64708 66660 64710
rect 66716 64708 66740 64710
rect 66796 64708 66820 64710
rect 66876 64708 66882 64710
rect 66574 64699 66882 64708
rect 5794 64220 6102 64229
rect 5794 64218 5800 64220
rect 5856 64218 5880 64220
rect 5936 64218 5960 64220
rect 6016 64218 6040 64220
rect 6096 64218 6102 64220
rect 5856 64166 5858 64218
rect 6038 64166 6040 64218
rect 5794 64164 5800 64166
rect 5856 64164 5880 64166
rect 5936 64164 5960 64166
rect 6016 64164 6040 64166
rect 6096 64164 6102 64166
rect 5794 64155 6102 64164
rect 36514 64220 36822 64229
rect 36514 64218 36520 64220
rect 36576 64218 36600 64220
rect 36656 64218 36680 64220
rect 36736 64218 36760 64220
rect 36816 64218 36822 64220
rect 36576 64166 36578 64218
rect 36758 64166 36760 64218
rect 36514 64164 36520 64166
rect 36576 64164 36600 64166
rect 36656 64164 36680 64166
rect 36736 64164 36760 64166
rect 36816 64164 36822 64166
rect 36514 64155 36822 64164
rect 67234 64220 67542 64229
rect 67234 64218 67240 64220
rect 67296 64218 67320 64220
rect 67376 64218 67400 64220
rect 67456 64218 67480 64220
rect 67536 64218 67542 64220
rect 67296 64166 67298 64218
rect 67478 64166 67480 64218
rect 67234 64164 67240 64166
rect 67296 64164 67320 64166
rect 67376 64164 67400 64166
rect 67456 64164 67480 64166
rect 67536 64164 67542 64166
rect 67234 64155 67542 64164
rect 5134 63676 5442 63685
rect 5134 63674 5140 63676
rect 5196 63674 5220 63676
rect 5276 63674 5300 63676
rect 5356 63674 5380 63676
rect 5436 63674 5442 63676
rect 5196 63622 5198 63674
rect 5378 63622 5380 63674
rect 5134 63620 5140 63622
rect 5196 63620 5220 63622
rect 5276 63620 5300 63622
rect 5356 63620 5380 63622
rect 5436 63620 5442 63622
rect 5134 63611 5442 63620
rect 35854 63676 36162 63685
rect 35854 63674 35860 63676
rect 35916 63674 35940 63676
rect 35996 63674 36020 63676
rect 36076 63674 36100 63676
rect 36156 63674 36162 63676
rect 35916 63622 35918 63674
rect 36098 63622 36100 63674
rect 35854 63620 35860 63622
rect 35916 63620 35940 63622
rect 35996 63620 36020 63622
rect 36076 63620 36100 63622
rect 36156 63620 36162 63622
rect 35854 63611 36162 63620
rect 66574 63676 66882 63685
rect 66574 63674 66580 63676
rect 66636 63674 66660 63676
rect 66716 63674 66740 63676
rect 66796 63674 66820 63676
rect 66876 63674 66882 63676
rect 66636 63622 66638 63674
rect 66818 63622 66820 63674
rect 66574 63620 66580 63622
rect 66636 63620 66660 63622
rect 66716 63620 66740 63622
rect 66796 63620 66820 63622
rect 66876 63620 66882 63622
rect 66574 63611 66882 63620
rect 5794 63132 6102 63141
rect 5794 63130 5800 63132
rect 5856 63130 5880 63132
rect 5936 63130 5960 63132
rect 6016 63130 6040 63132
rect 6096 63130 6102 63132
rect 5856 63078 5858 63130
rect 6038 63078 6040 63130
rect 5794 63076 5800 63078
rect 5856 63076 5880 63078
rect 5936 63076 5960 63078
rect 6016 63076 6040 63078
rect 6096 63076 6102 63078
rect 5794 63067 6102 63076
rect 36514 63132 36822 63141
rect 36514 63130 36520 63132
rect 36576 63130 36600 63132
rect 36656 63130 36680 63132
rect 36736 63130 36760 63132
rect 36816 63130 36822 63132
rect 36576 63078 36578 63130
rect 36758 63078 36760 63130
rect 36514 63076 36520 63078
rect 36576 63076 36600 63078
rect 36656 63076 36680 63078
rect 36736 63076 36760 63078
rect 36816 63076 36822 63078
rect 36514 63067 36822 63076
rect 67234 63132 67542 63141
rect 67234 63130 67240 63132
rect 67296 63130 67320 63132
rect 67376 63130 67400 63132
rect 67456 63130 67480 63132
rect 67536 63130 67542 63132
rect 67296 63078 67298 63130
rect 67478 63078 67480 63130
rect 67234 63076 67240 63078
rect 67296 63076 67320 63078
rect 67376 63076 67400 63078
rect 67456 63076 67480 63078
rect 67536 63076 67542 63078
rect 67234 63067 67542 63076
rect 5134 62588 5442 62597
rect 5134 62586 5140 62588
rect 5196 62586 5220 62588
rect 5276 62586 5300 62588
rect 5356 62586 5380 62588
rect 5436 62586 5442 62588
rect 5196 62534 5198 62586
rect 5378 62534 5380 62586
rect 5134 62532 5140 62534
rect 5196 62532 5220 62534
rect 5276 62532 5300 62534
rect 5356 62532 5380 62534
rect 5436 62532 5442 62534
rect 5134 62523 5442 62532
rect 35854 62588 36162 62597
rect 35854 62586 35860 62588
rect 35916 62586 35940 62588
rect 35996 62586 36020 62588
rect 36076 62586 36100 62588
rect 36156 62586 36162 62588
rect 35916 62534 35918 62586
rect 36098 62534 36100 62586
rect 35854 62532 35860 62534
rect 35916 62532 35940 62534
rect 35996 62532 36020 62534
rect 36076 62532 36100 62534
rect 36156 62532 36162 62534
rect 35854 62523 36162 62532
rect 66574 62588 66882 62597
rect 66574 62586 66580 62588
rect 66636 62586 66660 62588
rect 66716 62586 66740 62588
rect 66796 62586 66820 62588
rect 66876 62586 66882 62588
rect 66636 62534 66638 62586
rect 66818 62534 66820 62586
rect 66574 62532 66580 62534
rect 66636 62532 66660 62534
rect 66716 62532 66740 62534
rect 66796 62532 66820 62534
rect 66876 62532 66882 62534
rect 66574 62523 66882 62532
rect 5794 62044 6102 62053
rect 5794 62042 5800 62044
rect 5856 62042 5880 62044
rect 5936 62042 5960 62044
rect 6016 62042 6040 62044
rect 6096 62042 6102 62044
rect 5856 61990 5858 62042
rect 6038 61990 6040 62042
rect 5794 61988 5800 61990
rect 5856 61988 5880 61990
rect 5936 61988 5960 61990
rect 6016 61988 6040 61990
rect 6096 61988 6102 61990
rect 5794 61979 6102 61988
rect 36514 62044 36822 62053
rect 36514 62042 36520 62044
rect 36576 62042 36600 62044
rect 36656 62042 36680 62044
rect 36736 62042 36760 62044
rect 36816 62042 36822 62044
rect 36576 61990 36578 62042
rect 36758 61990 36760 62042
rect 36514 61988 36520 61990
rect 36576 61988 36600 61990
rect 36656 61988 36680 61990
rect 36736 61988 36760 61990
rect 36816 61988 36822 61990
rect 36514 61979 36822 61988
rect 67234 62044 67542 62053
rect 67234 62042 67240 62044
rect 67296 62042 67320 62044
rect 67376 62042 67400 62044
rect 67456 62042 67480 62044
rect 67536 62042 67542 62044
rect 67296 61990 67298 62042
rect 67478 61990 67480 62042
rect 67234 61988 67240 61990
rect 67296 61988 67320 61990
rect 67376 61988 67400 61990
rect 67456 61988 67480 61990
rect 67536 61988 67542 61990
rect 67234 61979 67542 61988
rect 5134 61500 5442 61509
rect 5134 61498 5140 61500
rect 5196 61498 5220 61500
rect 5276 61498 5300 61500
rect 5356 61498 5380 61500
rect 5436 61498 5442 61500
rect 5196 61446 5198 61498
rect 5378 61446 5380 61498
rect 5134 61444 5140 61446
rect 5196 61444 5220 61446
rect 5276 61444 5300 61446
rect 5356 61444 5380 61446
rect 5436 61444 5442 61446
rect 5134 61435 5442 61444
rect 35854 61500 36162 61509
rect 35854 61498 35860 61500
rect 35916 61498 35940 61500
rect 35996 61498 36020 61500
rect 36076 61498 36100 61500
rect 36156 61498 36162 61500
rect 35916 61446 35918 61498
rect 36098 61446 36100 61498
rect 35854 61444 35860 61446
rect 35916 61444 35940 61446
rect 35996 61444 36020 61446
rect 36076 61444 36100 61446
rect 36156 61444 36162 61446
rect 35854 61435 36162 61444
rect 66574 61500 66882 61509
rect 66574 61498 66580 61500
rect 66636 61498 66660 61500
rect 66716 61498 66740 61500
rect 66796 61498 66820 61500
rect 66876 61498 66882 61500
rect 66636 61446 66638 61498
rect 66818 61446 66820 61498
rect 66574 61444 66580 61446
rect 66636 61444 66660 61446
rect 66716 61444 66740 61446
rect 66796 61444 66820 61446
rect 66876 61444 66882 61446
rect 66574 61435 66882 61444
rect 5794 60956 6102 60965
rect 5794 60954 5800 60956
rect 5856 60954 5880 60956
rect 5936 60954 5960 60956
rect 6016 60954 6040 60956
rect 6096 60954 6102 60956
rect 5856 60902 5858 60954
rect 6038 60902 6040 60954
rect 5794 60900 5800 60902
rect 5856 60900 5880 60902
rect 5936 60900 5960 60902
rect 6016 60900 6040 60902
rect 6096 60900 6102 60902
rect 5794 60891 6102 60900
rect 36514 60956 36822 60965
rect 36514 60954 36520 60956
rect 36576 60954 36600 60956
rect 36656 60954 36680 60956
rect 36736 60954 36760 60956
rect 36816 60954 36822 60956
rect 36576 60902 36578 60954
rect 36758 60902 36760 60954
rect 36514 60900 36520 60902
rect 36576 60900 36600 60902
rect 36656 60900 36680 60902
rect 36736 60900 36760 60902
rect 36816 60900 36822 60902
rect 36514 60891 36822 60900
rect 67234 60956 67542 60965
rect 67234 60954 67240 60956
rect 67296 60954 67320 60956
rect 67376 60954 67400 60956
rect 67456 60954 67480 60956
rect 67536 60954 67542 60956
rect 67296 60902 67298 60954
rect 67478 60902 67480 60954
rect 67234 60900 67240 60902
rect 67296 60900 67320 60902
rect 67376 60900 67400 60902
rect 67456 60900 67480 60902
rect 67536 60900 67542 60902
rect 67234 60891 67542 60900
rect 5134 60412 5442 60421
rect 5134 60410 5140 60412
rect 5196 60410 5220 60412
rect 5276 60410 5300 60412
rect 5356 60410 5380 60412
rect 5436 60410 5442 60412
rect 5196 60358 5198 60410
rect 5378 60358 5380 60410
rect 5134 60356 5140 60358
rect 5196 60356 5220 60358
rect 5276 60356 5300 60358
rect 5356 60356 5380 60358
rect 5436 60356 5442 60358
rect 5134 60347 5442 60356
rect 35854 60412 36162 60421
rect 35854 60410 35860 60412
rect 35916 60410 35940 60412
rect 35996 60410 36020 60412
rect 36076 60410 36100 60412
rect 36156 60410 36162 60412
rect 35916 60358 35918 60410
rect 36098 60358 36100 60410
rect 35854 60356 35860 60358
rect 35916 60356 35940 60358
rect 35996 60356 36020 60358
rect 36076 60356 36100 60358
rect 36156 60356 36162 60358
rect 35854 60347 36162 60356
rect 66574 60412 66882 60421
rect 66574 60410 66580 60412
rect 66636 60410 66660 60412
rect 66716 60410 66740 60412
rect 66796 60410 66820 60412
rect 66876 60410 66882 60412
rect 66636 60358 66638 60410
rect 66818 60358 66820 60410
rect 66574 60356 66580 60358
rect 66636 60356 66660 60358
rect 66716 60356 66740 60358
rect 66796 60356 66820 60358
rect 66876 60356 66882 60358
rect 66574 60347 66882 60356
rect 5794 59868 6102 59877
rect 5794 59866 5800 59868
rect 5856 59866 5880 59868
rect 5936 59866 5960 59868
rect 6016 59866 6040 59868
rect 6096 59866 6102 59868
rect 5856 59814 5858 59866
rect 6038 59814 6040 59866
rect 5794 59812 5800 59814
rect 5856 59812 5880 59814
rect 5936 59812 5960 59814
rect 6016 59812 6040 59814
rect 6096 59812 6102 59814
rect 5794 59803 6102 59812
rect 36514 59868 36822 59877
rect 36514 59866 36520 59868
rect 36576 59866 36600 59868
rect 36656 59866 36680 59868
rect 36736 59866 36760 59868
rect 36816 59866 36822 59868
rect 36576 59814 36578 59866
rect 36758 59814 36760 59866
rect 36514 59812 36520 59814
rect 36576 59812 36600 59814
rect 36656 59812 36680 59814
rect 36736 59812 36760 59814
rect 36816 59812 36822 59814
rect 36514 59803 36822 59812
rect 67234 59868 67542 59877
rect 67234 59866 67240 59868
rect 67296 59866 67320 59868
rect 67376 59866 67400 59868
rect 67456 59866 67480 59868
rect 67536 59866 67542 59868
rect 67296 59814 67298 59866
rect 67478 59814 67480 59866
rect 67234 59812 67240 59814
rect 67296 59812 67320 59814
rect 67376 59812 67400 59814
rect 67456 59812 67480 59814
rect 67536 59812 67542 59814
rect 67234 59803 67542 59812
rect 5134 59324 5442 59333
rect 5134 59322 5140 59324
rect 5196 59322 5220 59324
rect 5276 59322 5300 59324
rect 5356 59322 5380 59324
rect 5436 59322 5442 59324
rect 5196 59270 5198 59322
rect 5378 59270 5380 59322
rect 5134 59268 5140 59270
rect 5196 59268 5220 59270
rect 5276 59268 5300 59270
rect 5356 59268 5380 59270
rect 5436 59268 5442 59270
rect 5134 59259 5442 59268
rect 35854 59324 36162 59333
rect 35854 59322 35860 59324
rect 35916 59322 35940 59324
rect 35996 59322 36020 59324
rect 36076 59322 36100 59324
rect 36156 59322 36162 59324
rect 35916 59270 35918 59322
rect 36098 59270 36100 59322
rect 35854 59268 35860 59270
rect 35916 59268 35940 59270
rect 35996 59268 36020 59270
rect 36076 59268 36100 59270
rect 36156 59268 36162 59270
rect 35854 59259 36162 59268
rect 66574 59324 66882 59333
rect 66574 59322 66580 59324
rect 66636 59322 66660 59324
rect 66716 59322 66740 59324
rect 66796 59322 66820 59324
rect 66876 59322 66882 59324
rect 66636 59270 66638 59322
rect 66818 59270 66820 59322
rect 66574 59268 66580 59270
rect 66636 59268 66660 59270
rect 66716 59268 66740 59270
rect 66796 59268 66820 59270
rect 66876 59268 66882 59270
rect 66574 59259 66882 59268
rect 5794 58780 6102 58789
rect 5794 58778 5800 58780
rect 5856 58778 5880 58780
rect 5936 58778 5960 58780
rect 6016 58778 6040 58780
rect 6096 58778 6102 58780
rect 5856 58726 5858 58778
rect 6038 58726 6040 58778
rect 5794 58724 5800 58726
rect 5856 58724 5880 58726
rect 5936 58724 5960 58726
rect 6016 58724 6040 58726
rect 6096 58724 6102 58726
rect 5794 58715 6102 58724
rect 36514 58780 36822 58789
rect 36514 58778 36520 58780
rect 36576 58778 36600 58780
rect 36656 58778 36680 58780
rect 36736 58778 36760 58780
rect 36816 58778 36822 58780
rect 36576 58726 36578 58778
rect 36758 58726 36760 58778
rect 36514 58724 36520 58726
rect 36576 58724 36600 58726
rect 36656 58724 36680 58726
rect 36736 58724 36760 58726
rect 36816 58724 36822 58726
rect 36514 58715 36822 58724
rect 67234 58780 67542 58789
rect 67234 58778 67240 58780
rect 67296 58778 67320 58780
rect 67376 58778 67400 58780
rect 67456 58778 67480 58780
rect 67536 58778 67542 58780
rect 67296 58726 67298 58778
rect 67478 58726 67480 58778
rect 67234 58724 67240 58726
rect 67296 58724 67320 58726
rect 67376 58724 67400 58726
rect 67456 58724 67480 58726
rect 67536 58724 67542 58726
rect 67234 58715 67542 58724
rect 5134 58236 5442 58245
rect 5134 58234 5140 58236
rect 5196 58234 5220 58236
rect 5276 58234 5300 58236
rect 5356 58234 5380 58236
rect 5436 58234 5442 58236
rect 5196 58182 5198 58234
rect 5378 58182 5380 58234
rect 5134 58180 5140 58182
rect 5196 58180 5220 58182
rect 5276 58180 5300 58182
rect 5356 58180 5380 58182
rect 5436 58180 5442 58182
rect 5134 58171 5442 58180
rect 35854 58236 36162 58245
rect 35854 58234 35860 58236
rect 35916 58234 35940 58236
rect 35996 58234 36020 58236
rect 36076 58234 36100 58236
rect 36156 58234 36162 58236
rect 35916 58182 35918 58234
rect 36098 58182 36100 58234
rect 35854 58180 35860 58182
rect 35916 58180 35940 58182
rect 35996 58180 36020 58182
rect 36076 58180 36100 58182
rect 36156 58180 36162 58182
rect 35854 58171 36162 58180
rect 66574 58236 66882 58245
rect 66574 58234 66580 58236
rect 66636 58234 66660 58236
rect 66716 58234 66740 58236
rect 66796 58234 66820 58236
rect 66876 58234 66882 58236
rect 66636 58182 66638 58234
rect 66818 58182 66820 58234
rect 66574 58180 66580 58182
rect 66636 58180 66660 58182
rect 66716 58180 66740 58182
rect 66796 58180 66820 58182
rect 66876 58180 66882 58182
rect 66574 58171 66882 58180
rect 5794 57692 6102 57701
rect 5794 57690 5800 57692
rect 5856 57690 5880 57692
rect 5936 57690 5960 57692
rect 6016 57690 6040 57692
rect 6096 57690 6102 57692
rect 5856 57638 5858 57690
rect 6038 57638 6040 57690
rect 5794 57636 5800 57638
rect 5856 57636 5880 57638
rect 5936 57636 5960 57638
rect 6016 57636 6040 57638
rect 6096 57636 6102 57638
rect 5794 57627 6102 57636
rect 36514 57692 36822 57701
rect 36514 57690 36520 57692
rect 36576 57690 36600 57692
rect 36656 57690 36680 57692
rect 36736 57690 36760 57692
rect 36816 57690 36822 57692
rect 36576 57638 36578 57690
rect 36758 57638 36760 57690
rect 36514 57636 36520 57638
rect 36576 57636 36600 57638
rect 36656 57636 36680 57638
rect 36736 57636 36760 57638
rect 36816 57636 36822 57638
rect 36514 57627 36822 57636
rect 67234 57692 67542 57701
rect 67234 57690 67240 57692
rect 67296 57690 67320 57692
rect 67376 57690 67400 57692
rect 67456 57690 67480 57692
rect 67536 57690 67542 57692
rect 67296 57638 67298 57690
rect 67478 57638 67480 57690
rect 67234 57636 67240 57638
rect 67296 57636 67320 57638
rect 67376 57636 67400 57638
rect 67456 57636 67480 57638
rect 67536 57636 67542 57638
rect 67234 57627 67542 57636
rect 5134 57148 5442 57157
rect 5134 57146 5140 57148
rect 5196 57146 5220 57148
rect 5276 57146 5300 57148
rect 5356 57146 5380 57148
rect 5436 57146 5442 57148
rect 5196 57094 5198 57146
rect 5378 57094 5380 57146
rect 5134 57092 5140 57094
rect 5196 57092 5220 57094
rect 5276 57092 5300 57094
rect 5356 57092 5380 57094
rect 5436 57092 5442 57094
rect 5134 57083 5442 57092
rect 35854 57148 36162 57157
rect 35854 57146 35860 57148
rect 35916 57146 35940 57148
rect 35996 57146 36020 57148
rect 36076 57146 36100 57148
rect 36156 57146 36162 57148
rect 35916 57094 35918 57146
rect 36098 57094 36100 57146
rect 35854 57092 35860 57094
rect 35916 57092 35940 57094
rect 35996 57092 36020 57094
rect 36076 57092 36100 57094
rect 36156 57092 36162 57094
rect 35854 57083 36162 57092
rect 66574 57148 66882 57157
rect 66574 57146 66580 57148
rect 66636 57146 66660 57148
rect 66716 57146 66740 57148
rect 66796 57146 66820 57148
rect 66876 57146 66882 57148
rect 66636 57094 66638 57146
rect 66818 57094 66820 57146
rect 66574 57092 66580 57094
rect 66636 57092 66660 57094
rect 66716 57092 66740 57094
rect 66796 57092 66820 57094
rect 66876 57092 66882 57094
rect 66574 57083 66882 57092
rect 5794 56604 6102 56613
rect 5794 56602 5800 56604
rect 5856 56602 5880 56604
rect 5936 56602 5960 56604
rect 6016 56602 6040 56604
rect 6096 56602 6102 56604
rect 5856 56550 5858 56602
rect 6038 56550 6040 56602
rect 5794 56548 5800 56550
rect 5856 56548 5880 56550
rect 5936 56548 5960 56550
rect 6016 56548 6040 56550
rect 6096 56548 6102 56550
rect 5794 56539 6102 56548
rect 36514 56604 36822 56613
rect 36514 56602 36520 56604
rect 36576 56602 36600 56604
rect 36656 56602 36680 56604
rect 36736 56602 36760 56604
rect 36816 56602 36822 56604
rect 36576 56550 36578 56602
rect 36758 56550 36760 56602
rect 36514 56548 36520 56550
rect 36576 56548 36600 56550
rect 36656 56548 36680 56550
rect 36736 56548 36760 56550
rect 36816 56548 36822 56550
rect 36514 56539 36822 56548
rect 67234 56604 67542 56613
rect 67234 56602 67240 56604
rect 67296 56602 67320 56604
rect 67376 56602 67400 56604
rect 67456 56602 67480 56604
rect 67536 56602 67542 56604
rect 67296 56550 67298 56602
rect 67478 56550 67480 56602
rect 67234 56548 67240 56550
rect 67296 56548 67320 56550
rect 67376 56548 67400 56550
rect 67456 56548 67480 56550
rect 67536 56548 67542 56550
rect 67234 56539 67542 56548
rect 5134 56060 5442 56069
rect 5134 56058 5140 56060
rect 5196 56058 5220 56060
rect 5276 56058 5300 56060
rect 5356 56058 5380 56060
rect 5436 56058 5442 56060
rect 5196 56006 5198 56058
rect 5378 56006 5380 56058
rect 5134 56004 5140 56006
rect 5196 56004 5220 56006
rect 5276 56004 5300 56006
rect 5356 56004 5380 56006
rect 5436 56004 5442 56006
rect 5134 55995 5442 56004
rect 35854 56060 36162 56069
rect 35854 56058 35860 56060
rect 35916 56058 35940 56060
rect 35996 56058 36020 56060
rect 36076 56058 36100 56060
rect 36156 56058 36162 56060
rect 35916 56006 35918 56058
rect 36098 56006 36100 56058
rect 35854 56004 35860 56006
rect 35916 56004 35940 56006
rect 35996 56004 36020 56006
rect 36076 56004 36100 56006
rect 36156 56004 36162 56006
rect 35854 55995 36162 56004
rect 66574 56060 66882 56069
rect 66574 56058 66580 56060
rect 66636 56058 66660 56060
rect 66716 56058 66740 56060
rect 66796 56058 66820 56060
rect 66876 56058 66882 56060
rect 66636 56006 66638 56058
rect 66818 56006 66820 56058
rect 66574 56004 66580 56006
rect 66636 56004 66660 56006
rect 66716 56004 66740 56006
rect 66796 56004 66820 56006
rect 66876 56004 66882 56006
rect 66574 55995 66882 56004
rect 5794 55516 6102 55525
rect 5794 55514 5800 55516
rect 5856 55514 5880 55516
rect 5936 55514 5960 55516
rect 6016 55514 6040 55516
rect 6096 55514 6102 55516
rect 5856 55462 5858 55514
rect 6038 55462 6040 55514
rect 5794 55460 5800 55462
rect 5856 55460 5880 55462
rect 5936 55460 5960 55462
rect 6016 55460 6040 55462
rect 6096 55460 6102 55462
rect 5794 55451 6102 55460
rect 36514 55516 36822 55525
rect 36514 55514 36520 55516
rect 36576 55514 36600 55516
rect 36656 55514 36680 55516
rect 36736 55514 36760 55516
rect 36816 55514 36822 55516
rect 36576 55462 36578 55514
rect 36758 55462 36760 55514
rect 36514 55460 36520 55462
rect 36576 55460 36600 55462
rect 36656 55460 36680 55462
rect 36736 55460 36760 55462
rect 36816 55460 36822 55462
rect 36514 55451 36822 55460
rect 67234 55516 67542 55525
rect 67234 55514 67240 55516
rect 67296 55514 67320 55516
rect 67376 55514 67400 55516
rect 67456 55514 67480 55516
rect 67536 55514 67542 55516
rect 67296 55462 67298 55514
rect 67478 55462 67480 55514
rect 67234 55460 67240 55462
rect 67296 55460 67320 55462
rect 67376 55460 67400 55462
rect 67456 55460 67480 55462
rect 67536 55460 67542 55462
rect 67234 55451 67542 55460
rect 5134 54972 5442 54981
rect 5134 54970 5140 54972
rect 5196 54970 5220 54972
rect 5276 54970 5300 54972
rect 5356 54970 5380 54972
rect 5436 54970 5442 54972
rect 5196 54918 5198 54970
rect 5378 54918 5380 54970
rect 5134 54916 5140 54918
rect 5196 54916 5220 54918
rect 5276 54916 5300 54918
rect 5356 54916 5380 54918
rect 5436 54916 5442 54918
rect 5134 54907 5442 54916
rect 35854 54972 36162 54981
rect 35854 54970 35860 54972
rect 35916 54970 35940 54972
rect 35996 54970 36020 54972
rect 36076 54970 36100 54972
rect 36156 54970 36162 54972
rect 35916 54918 35918 54970
rect 36098 54918 36100 54970
rect 35854 54916 35860 54918
rect 35916 54916 35940 54918
rect 35996 54916 36020 54918
rect 36076 54916 36100 54918
rect 36156 54916 36162 54918
rect 35854 54907 36162 54916
rect 66574 54972 66882 54981
rect 66574 54970 66580 54972
rect 66636 54970 66660 54972
rect 66716 54970 66740 54972
rect 66796 54970 66820 54972
rect 66876 54970 66882 54972
rect 66636 54918 66638 54970
rect 66818 54918 66820 54970
rect 66574 54916 66580 54918
rect 66636 54916 66660 54918
rect 66716 54916 66740 54918
rect 66796 54916 66820 54918
rect 66876 54916 66882 54918
rect 66574 54907 66882 54916
rect 5794 54428 6102 54437
rect 5794 54426 5800 54428
rect 5856 54426 5880 54428
rect 5936 54426 5960 54428
rect 6016 54426 6040 54428
rect 6096 54426 6102 54428
rect 5856 54374 5858 54426
rect 6038 54374 6040 54426
rect 5794 54372 5800 54374
rect 5856 54372 5880 54374
rect 5936 54372 5960 54374
rect 6016 54372 6040 54374
rect 6096 54372 6102 54374
rect 5794 54363 6102 54372
rect 36514 54428 36822 54437
rect 36514 54426 36520 54428
rect 36576 54426 36600 54428
rect 36656 54426 36680 54428
rect 36736 54426 36760 54428
rect 36816 54426 36822 54428
rect 36576 54374 36578 54426
rect 36758 54374 36760 54426
rect 36514 54372 36520 54374
rect 36576 54372 36600 54374
rect 36656 54372 36680 54374
rect 36736 54372 36760 54374
rect 36816 54372 36822 54374
rect 36514 54363 36822 54372
rect 67234 54428 67542 54437
rect 67234 54426 67240 54428
rect 67296 54426 67320 54428
rect 67376 54426 67400 54428
rect 67456 54426 67480 54428
rect 67536 54426 67542 54428
rect 67296 54374 67298 54426
rect 67478 54374 67480 54426
rect 67234 54372 67240 54374
rect 67296 54372 67320 54374
rect 67376 54372 67400 54374
rect 67456 54372 67480 54374
rect 67536 54372 67542 54374
rect 67234 54363 67542 54372
rect 5134 53884 5442 53893
rect 5134 53882 5140 53884
rect 5196 53882 5220 53884
rect 5276 53882 5300 53884
rect 5356 53882 5380 53884
rect 5436 53882 5442 53884
rect 5196 53830 5198 53882
rect 5378 53830 5380 53882
rect 5134 53828 5140 53830
rect 5196 53828 5220 53830
rect 5276 53828 5300 53830
rect 5356 53828 5380 53830
rect 5436 53828 5442 53830
rect 5134 53819 5442 53828
rect 35854 53884 36162 53893
rect 35854 53882 35860 53884
rect 35916 53882 35940 53884
rect 35996 53882 36020 53884
rect 36076 53882 36100 53884
rect 36156 53882 36162 53884
rect 35916 53830 35918 53882
rect 36098 53830 36100 53882
rect 35854 53828 35860 53830
rect 35916 53828 35940 53830
rect 35996 53828 36020 53830
rect 36076 53828 36100 53830
rect 36156 53828 36162 53830
rect 35854 53819 36162 53828
rect 66574 53884 66882 53893
rect 66574 53882 66580 53884
rect 66636 53882 66660 53884
rect 66716 53882 66740 53884
rect 66796 53882 66820 53884
rect 66876 53882 66882 53884
rect 66636 53830 66638 53882
rect 66818 53830 66820 53882
rect 66574 53828 66580 53830
rect 66636 53828 66660 53830
rect 66716 53828 66740 53830
rect 66796 53828 66820 53830
rect 66876 53828 66882 53830
rect 66574 53819 66882 53828
rect 5794 53340 6102 53349
rect 5794 53338 5800 53340
rect 5856 53338 5880 53340
rect 5936 53338 5960 53340
rect 6016 53338 6040 53340
rect 6096 53338 6102 53340
rect 5856 53286 5858 53338
rect 6038 53286 6040 53338
rect 5794 53284 5800 53286
rect 5856 53284 5880 53286
rect 5936 53284 5960 53286
rect 6016 53284 6040 53286
rect 6096 53284 6102 53286
rect 5794 53275 6102 53284
rect 36514 53340 36822 53349
rect 36514 53338 36520 53340
rect 36576 53338 36600 53340
rect 36656 53338 36680 53340
rect 36736 53338 36760 53340
rect 36816 53338 36822 53340
rect 36576 53286 36578 53338
rect 36758 53286 36760 53338
rect 36514 53284 36520 53286
rect 36576 53284 36600 53286
rect 36656 53284 36680 53286
rect 36736 53284 36760 53286
rect 36816 53284 36822 53286
rect 36514 53275 36822 53284
rect 67234 53340 67542 53349
rect 67234 53338 67240 53340
rect 67296 53338 67320 53340
rect 67376 53338 67400 53340
rect 67456 53338 67480 53340
rect 67536 53338 67542 53340
rect 67296 53286 67298 53338
rect 67478 53286 67480 53338
rect 67234 53284 67240 53286
rect 67296 53284 67320 53286
rect 67376 53284 67400 53286
rect 67456 53284 67480 53286
rect 67536 53284 67542 53286
rect 67234 53275 67542 53284
rect 5134 52796 5442 52805
rect 5134 52794 5140 52796
rect 5196 52794 5220 52796
rect 5276 52794 5300 52796
rect 5356 52794 5380 52796
rect 5436 52794 5442 52796
rect 5196 52742 5198 52794
rect 5378 52742 5380 52794
rect 5134 52740 5140 52742
rect 5196 52740 5220 52742
rect 5276 52740 5300 52742
rect 5356 52740 5380 52742
rect 5436 52740 5442 52742
rect 5134 52731 5442 52740
rect 35854 52796 36162 52805
rect 35854 52794 35860 52796
rect 35916 52794 35940 52796
rect 35996 52794 36020 52796
rect 36076 52794 36100 52796
rect 36156 52794 36162 52796
rect 35916 52742 35918 52794
rect 36098 52742 36100 52794
rect 35854 52740 35860 52742
rect 35916 52740 35940 52742
rect 35996 52740 36020 52742
rect 36076 52740 36100 52742
rect 36156 52740 36162 52742
rect 35854 52731 36162 52740
rect 66574 52796 66882 52805
rect 66574 52794 66580 52796
rect 66636 52794 66660 52796
rect 66716 52794 66740 52796
rect 66796 52794 66820 52796
rect 66876 52794 66882 52796
rect 66636 52742 66638 52794
rect 66818 52742 66820 52794
rect 66574 52740 66580 52742
rect 66636 52740 66660 52742
rect 66716 52740 66740 52742
rect 66796 52740 66820 52742
rect 66876 52740 66882 52742
rect 66574 52731 66882 52740
rect 5794 52252 6102 52261
rect 5794 52250 5800 52252
rect 5856 52250 5880 52252
rect 5936 52250 5960 52252
rect 6016 52250 6040 52252
rect 6096 52250 6102 52252
rect 5856 52198 5858 52250
rect 6038 52198 6040 52250
rect 5794 52196 5800 52198
rect 5856 52196 5880 52198
rect 5936 52196 5960 52198
rect 6016 52196 6040 52198
rect 6096 52196 6102 52198
rect 5794 52187 6102 52196
rect 36514 52252 36822 52261
rect 36514 52250 36520 52252
rect 36576 52250 36600 52252
rect 36656 52250 36680 52252
rect 36736 52250 36760 52252
rect 36816 52250 36822 52252
rect 36576 52198 36578 52250
rect 36758 52198 36760 52250
rect 36514 52196 36520 52198
rect 36576 52196 36600 52198
rect 36656 52196 36680 52198
rect 36736 52196 36760 52198
rect 36816 52196 36822 52198
rect 36514 52187 36822 52196
rect 67234 52252 67542 52261
rect 67234 52250 67240 52252
rect 67296 52250 67320 52252
rect 67376 52250 67400 52252
rect 67456 52250 67480 52252
rect 67536 52250 67542 52252
rect 67296 52198 67298 52250
rect 67478 52198 67480 52250
rect 67234 52196 67240 52198
rect 67296 52196 67320 52198
rect 67376 52196 67400 52198
rect 67456 52196 67480 52198
rect 67536 52196 67542 52198
rect 67234 52187 67542 52196
rect 77576 51808 77628 51814
rect 77574 51776 77576 51785
rect 77628 51776 77630 51785
rect 5134 51708 5442 51717
rect 5134 51706 5140 51708
rect 5196 51706 5220 51708
rect 5276 51706 5300 51708
rect 5356 51706 5380 51708
rect 5436 51706 5442 51708
rect 5196 51654 5198 51706
rect 5378 51654 5380 51706
rect 5134 51652 5140 51654
rect 5196 51652 5220 51654
rect 5276 51652 5300 51654
rect 5356 51652 5380 51654
rect 5436 51652 5442 51654
rect 5134 51643 5442 51652
rect 35854 51708 36162 51717
rect 35854 51706 35860 51708
rect 35916 51706 35940 51708
rect 35996 51706 36020 51708
rect 36076 51706 36100 51708
rect 36156 51706 36162 51708
rect 35916 51654 35918 51706
rect 36098 51654 36100 51706
rect 35854 51652 35860 51654
rect 35916 51652 35940 51654
rect 35996 51652 36020 51654
rect 36076 51652 36100 51654
rect 36156 51652 36162 51654
rect 35854 51643 36162 51652
rect 66574 51708 66882 51717
rect 77574 51711 77630 51720
rect 66574 51706 66580 51708
rect 66636 51706 66660 51708
rect 66716 51706 66740 51708
rect 66796 51706 66820 51708
rect 66876 51706 66882 51708
rect 66636 51654 66638 51706
rect 66818 51654 66820 51706
rect 66574 51652 66580 51654
rect 66636 51652 66660 51654
rect 66716 51652 66740 51654
rect 66796 51652 66820 51654
rect 66876 51652 66882 51654
rect 66574 51643 66882 51652
rect 5794 51164 6102 51173
rect 5794 51162 5800 51164
rect 5856 51162 5880 51164
rect 5936 51162 5960 51164
rect 6016 51162 6040 51164
rect 6096 51162 6102 51164
rect 5856 51110 5858 51162
rect 6038 51110 6040 51162
rect 5794 51108 5800 51110
rect 5856 51108 5880 51110
rect 5936 51108 5960 51110
rect 6016 51108 6040 51110
rect 6096 51108 6102 51110
rect 5794 51099 6102 51108
rect 36514 51164 36822 51173
rect 36514 51162 36520 51164
rect 36576 51162 36600 51164
rect 36656 51162 36680 51164
rect 36736 51162 36760 51164
rect 36816 51162 36822 51164
rect 36576 51110 36578 51162
rect 36758 51110 36760 51162
rect 36514 51108 36520 51110
rect 36576 51108 36600 51110
rect 36656 51108 36680 51110
rect 36736 51108 36760 51110
rect 36816 51108 36822 51110
rect 36514 51099 36822 51108
rect 67234 51164 67542 51173
rect 67234 51162 67240 51164
rect 67296 51162 67320 51164
rect 67376 51162 67400 51164
rect 67456 51162 67480 51164
rect 67536 51162 67542 51164
rect 67296 51110 67298 51162
rect 67478 51110 67480 51162
rect 67234 51108 67240 51110
rect 67296 51108 67320 51110
rect 67376 51108 67400 51110
rect 67456 51108 67480 51110
rect 67536 51108 67542 51110
rect 67234 51099 67542 51108
rect 5134 50620 5442 50629
rect 5134 50618 5140 50620
rect 5196 50618 5220 50620
rect 5276 50618 5300 50620
rect 5356 50618 5380 50620
rect 5436 50618 5442 50620
rect 5196 50566 5198 50618
rect 5378 50566 5380 50618
rect 5134 50564 5140 50566
rect 5196 50564 5220 50566
rect 5276 50564 5300 50566
rect 5356 50564 5380 50566
rect 5436 50564 5442 50566
rect 5134 50555 5442 50564
rect 35854 50620 36162 50629
rect 35854 50618 35860 50620
rect 35916 50618 35940 50620
rect 35996 50618 36020 50620
rect 36076 50618 36100 50620
rect 36156 50618 36162 50620
rect 35916 50566 35918 50618
rect 36098 50566 36100 50618
rect 35854 50564 35860 50566
rect 35916 50564 35940 50566
rect 35996 50564 36020 50566
rect 36076 50564 36100 50566
rect 36156 50564 36162 50566
rect 35854 50555 36162 50564
rect 66574 50620 66882 50629
rect 66574 50618 66580 50620
rect 66636 50618 66660 50620
rect 66716 50618 66740 50620
rect 66796 50618 66820 50620
rect 66876 50618 66882 50620
rect 66636 50566 66638 50618
rect 66818 50566 66820 50618
rect 66574 50564 66580 50566
rect 66636 50564 66660 50566
rect 66716 50564 66740 50566
rect 66796 50564 66820 50566
rect 66876 50564 66882 50566
rect 66574 50555 66882 50564
rect 5794 50076 6102 50085
rect 5794 50074 5800 50076
rect 5856 50074 5880 50076
rect 5936 50074 5960 50076
rect 6016 50074 6040 50076
rect 6096 50074 6102 50076
rect 5856 50022 5858 50074
rect 6038 50022 6040 50074
rect 5794 50020 5800 50022
rect 5856 50020 5880 50022
rect 5936 50020 5960 50022
rect 6016 50020 6040 50022
rect 6096 50020 6102 50022
rect 5794 50011 6102 50020
rect 36514 50076 36822 50085
rect 36514 50074 36520 50076
rect 36576 50074 36600 50076
rect 36656 50074 36680 50076
rect 36736 50074 36760 50076
rect 36816 50074 36822 50076
rect 36576 50022 36578 50074
rect 36758 50022 36760 50074
rect 36514 50020 36520 50022
rect 36576 50020 36600 50022
rect 36656 50020 36680 50022
rect 36736 50020 36760 50022
rect 36816 50020 36822 50022
rect 36514 50011 36822 50020
rect 67234 50076 67542 50085
rect 67234 50074 67240 50076
rect 67296 50074 67320 50076
rect 67376 50074 67400 50076
rect 67456 50074 67480 50076
rect 67536 50074 67542 50076
rect 67296 50022 67298 50074
rect 67478 50022 67480 50074
rect 67234 50020 67240 50022
rect 67296 50020 67320 50022
rect 67376 50020 67400 50022
rect 67456 50020 67480 50022
rect 67536 50020 67542 50022
rect 67234 50011 67542 50020
rect 77576 49768 77628 49774
rect 77574 49736 77576 49745
rect 77628 49736 77630 49745
rect 77574 49671 77630 49680
rect 5134 49532 5442 49541
rect 5134 49530 5140 49532
rect 5196 49530 5220 49532
rect 5276 49530 5300 49532
rect 5356 49530 5380 49532
rect 5436 49530 5442 49532
rect 5196 49478 5198 49530
rect 5378 49478 5380 49530
rect 5134 49476 5140 49478
rect 5196 49476 5220 49478
rect 5276 49476 5300 49478
rect 5356 49476 5380 49478
rect 5436 49476 5442 49478
rect 5134 49467 5442 49476
rect 35854 49532 36162 49541
rect 35854 49530 35860 49532
rect 35916 49530 35940 49532
rect 35996 49530 36020 49532
rect 36076 49530 36100 49532
rect 36156 49530 36162 49532
rect 35916 49478 35918 49530
rect 36098 49478 36100 49530
rect 35854 49476 35860 49478
rect 35916 49476 35940 49478
rect 35996 49476 36020 49478
rect 36076 49476 36100 49478
rect 36156 49476 36162 49478
rect 35854 49467 36162 49476
rect 66574 49532 66882 49541
rect 66574 49530 66580 49532
rect 66636 49530 66660 49532
rect 66716 49530 66740 49532
rect 66796 49530 66820 49532
rect 66876 49530 66882 49532
rect 66636 49478 66638 49530
rect 66818 49478 66820 49530
rect 66574 49476 66580 49478
rect 66636 49476 66660 49478
rect 66716 49476 66740 49478
rect 66796 49476 66820 49478
rect 66876 49476 66882 49478
rect 66574 49467 66882 49476
rect 5794 48988 6102 48997
rect 5794 48986 5800 48988
rect 5856 48986 5880 48988
rect 5936 48986 5960 48988
rect 6016 48986 6040 48988
rect 6096 48986 6102 48988
rect 5856 48934 5858 48986
rect 6038 48934 6040 48986
rect 5794 48932 5800 48934
rect 5856 48932 5880 48934
rect 5936 48932 5960 48934
rect 6016 48932 6040 48934
rect 6096 48932 6102 48934
rect 5794 48923 6102 48932
rect 36514 48988 36822 48997
rect 36514 48986 36520 48988
rect 36576 48986 36600 48988
rect 36656 48986 36680 48988
rect 36736 48986 36760 48988
rect 36816 48986 36822 48988
rect 36576 48934 36578 48986
rect 36758 48934 36760 48986
rect 36514 48932 36520 48934
rect 36576 48932 36600 48934
rect 36656 48932 36680 48934
rect 36736 48932 36760 48934
rect 36816 48932 36822 48934
rect 36514 48923 36822 48932
rect 67234 48988 67542 48997
rect 67234 48986 67240 48988
rect 67296 48986 67320 48988
rect 67376 48986 67400 48988
rect 67456 48986 67480 48988
rect 67536 48986 67542 48988
rect 67296 48934 67298 48986
rect 67478 48934 67480 48986
rect 67234 48932 67240 48934
rect 67296 48932 67320 48934
rect 67376 48932 67400 48934
rect 67456 48932 67480 48934
rect 67536 48932 67542 48934
rect 67234 48923 67542 48932
rect 5134 48444 5442 48453
rect 5134 48442 5140 48444
rect 5196 48442 5220 48444
rect 5276 48442 5300 48444
rect 5356 48442 5380 48444
rect 5436 48442 5442 48444
rect 5196 48390 5198 48442
rect 5378 48390 5380 48442
rect 5134 48388 5140 48390
rect 5196 48388 5220 48390
rect 5276 48388 5300 48390
rect 5356 48388 5380 48390
rect 5436 48388 5442 48390
rect 5134 48379 5442 48388
rect 35854 48444 36162 48453
rect 35854 48442 35860 48444
rect 35916 48442 35940 48444
rect 35996 48442 36020 48444
rect 36076 48442 36100 48444
rect 36156 48442 36162 48444
rect 35916 48390 35918 48442
rect 36098 48390 36100 48442
rect 35854 48388 35860 48390
rect 35916 48388 35940 48390
rect 35996 48388 36020 48390
rect 36076 48388 36100 48390
rect 36156 48388 36162 48390
rect 35854 48379 36162 48388
rect 66574 48444 66882 48453
rect 66574 48442 66580 48444
rect 66636 48442 66660 48444
rect 66716 48442 66740 48444
rect 66796 48442 66820 48444
rect 66876 48442 66882 48444
rect 66636 48390 66638 48442
rect 66818 48390 66820 48442
rect 66574 48388 66580 48390
rect 66636 48388 66660 48390
rect 66716 48388 66740 48390
rect 66796 48388 66820 48390
rect 66876 48388 66882 48390
rect 66574 48379 66882 48388
rect 5794 47900 6102 47909
rect 5794 47898 5800 47900
rect 5856 47898 5880 47900
rect 5936 47898 5960 47900
rect 6016 47898 6040 47900
rect 6096 47898 6102 47900
rect 5856 47846 5858 47898
rect 6038 47846 6040 47898
rect 5794 47844 5800 47846
rect 5856 47844 5880 47846
rect 5936 47844 5960 47846
rect 6016 47844 6040 47846
rect 6096 47844 6102 47846
rect 5794 47835 6102 47844
rect 36514 47900 36822 47909
rect 36514 47898 36520 47900
rect 36576 47898 36600 47900
rect 36656 47898 36680 47900
rect 36736 47898 36760 47900
rect 36816 47898 36822 47900
rect 36576 47846 36578 47898
rect 36758 47846 36760 47898
rect 36514 47844 36520 47846
rect 36576 47844 36600 47846
rect 36656 47844 36680 47846
rect 36736 47844 36760 47846
rect 36816 47844 36822 47846
rect 36514 47835 36822 47844
rect 67234 47900 67542 47909
rect 67234 47898 67240 47900
rect 67296 47898 67320 47900
rect 67376 47898 67400 47900
rect 67456 47898 67480 47900
rect 67536 47898 67542 47900
rect 67296 47846 67298 47898
rect 67478 47846 67480 47898
rect 67234 47844 67240 47846
rect 67296 47844 67320 47846
rect 67376 47844 67400 47846
rect 67456 47844 67480 47846
rect 67536 47844 67542 47846
rect 67234 47835 67542 47844
rect 5134 47356 5442 47365
rect 5134 47354 5140 47356
rect 5196 47354 5220 47356
rect 5276 47354 5300 47356
rect 5356 47354 5380 47356
rect 5436 47354 5442 47356
rect 5196 47302 5198 47354
rect 5378 47302 5380 47354
rect 5134 47300 5140 47302
rect 5196 47300 5220 47302
rect 5276 47300 5300 47302
rect 5356 47300 5380 47302
rect 5436 47300 5442 47302
rect 5134 47291 5442 47300
rect 35854 47356 36162 47365
rect 35854 47354 35860 47356
rect 35916 47354 35940 47356
rect 35996 47354 36020 47356
rect 36076 47354 36100 47356
rect 36156 47354 36162 47356
rect 35916 47302 35918 47354
rect 36098 47302 36100 47354
rect 35854 47300 35860 47302
rect 35916 47300 35940 47302
rect 35996 47300 36020 47302
rect 36076 47300 36100 47302
rect 36156 47300 36162 47302
rect 35854 47291 36162 47300
rect 66574 47356 66882 47365
rect 66574 47354 66580 47356
rect 66636 47354 66660 47356
rect 66716 47354 66740 47356
rect 66796 47354 66820 47356
rect 66876 47354 66882 47356
rect 66636 47302 66638 47354
rect 66818 47302 66820 47354
rect 66574 47300 66580 47302
rect 66636 47300 66660 47302
rect 66716 47300 66740 47302
rect 66796 47300 66820 47302
rect 66876 47300 66882 47302
rect 66574 47291 66882 47300
rect 5794 46812 6102 46821
rect 5794 46810 5800 46812
rect 5856 46810 5880 46812
rect 5936 46810 5960 46812
rect 6016 46810 6040 46812
rect 6096 46810 6102 46812
rect 5856 46758 5858 46810
rect 6038 46758 6040 46810
rect 5794 46756 5800 46758
rect 5856 46756 5880 46758
rect 5936 46756 5960 46758
rect 6016 46756 6040 46758
rect 6096 46756 6102 46758
rect 5794 46747 6102 46756
rect 36514 46812 36822 46821
rect 36514 46810 36520 46812
rect 36576 46810 36600 46812
rect 36656 46810 36680 46812
rect 36736 46810 36760 46812
rect 36816 46810 36822 46812
rect 36576 46758 36578 46810
rect 36758 46758 36760 46810
rect 36514 46756 36520 46758
rect 36576 46756 36600 46758
rect 36656 46756 36680 46758
rect 36736 46756 36760 46758
rect 36816 46756 36822 46758
rect 36514 46747 36822 46756
rect 67234 46812 67542 46821
rect 67234 46810 67240 46812
rect 67296 46810 67320 46812
rect 67376 46810 67400 46812
rect 67456 46810 67480 46812
rect 67536 46810 67542 46812
rect 67296 46758 67298 46810
rect 67478 46758 67480 46810
rect 67234 46756 67240 46758
rect 67296 46756 67320 46758
rect 67376 46756 67400 46758
rect 67456 46756 67480 46758
rect 67536 46756 67542 46758
rect 67234 46747 67542 46756
rect 5134 46268 5442 46277
rect 5134 46266 5140 46268
rect 5196 46266 5220 46268
rect 5276 46266 5300 46268
rect 5356 46266 5380 46268
rect 5436 46266 5442 46268
rect 5196 46214 5198 46266
rect 5378 46214 5380 46266
rect 5134 46212 5140 46214
rect 5196 46212 5220 46214
rect 5276 46212 5300 46214
rect 5356 46212 5380 46214
rect 5436 46212 5442 46214
rect 5134 46203 5442 46212
rect 35854 46268 36162 46277
rect 35854 46266 35860 46268
rect 35916 46266 35940 46268
rect 35996 46266 36020 46268
rect 36076 46266 36100 46268
rect 36156 46266 36162 46268
rect 35916 46214 35918 46266
rect 36098 46214 36100 46266
rect 35854 46212 35860 46214
rect 35916 46212 35940 46214
rect 35996 46212 36020 46214
rect 36076 46212 36100 46214
rect 36156 46212 36162 46214
rect 35854 46203 36162 46212
rect 66574 46268 66882 46277
rect 66574 46266 66580 46268
rect 66636 46266 66660 46268
rect 66716 46266 66740 46268
rect 66796 46266 66820 46268
rect 66876 46266 66882 46268
rect 66636 46214 66638 46266
rect 66818 46214 66820 46266
rect 66574 46212 66580 46214
rect 66636 46212 66660 46214
rect 66716 46212 66740 46214
rect 66796 46212 66820 46214
rect 66876 46212 66882 46214
rect 66574 46203 66882 46212
rect 5794 45724 6102 45733
rect 5794 45722 5800 45724
rect 5856 45722 5880 45724
rect 5936 45722 5960 45724
rect 6016 45722 6040 45724
rect 6096 45722 6102 45724
rect 5856 45670 5858 45722
rect 6038 45670 6040 45722
rect 5794 45668 5800 45670
rect 5856 45668 5880 45670
rect 5936 45668 5960 45670
rect 6016 45668 6040 45670
rect 6096 45668 6102 45670
rect 1306 45656 1362 45665
rect 5794 45659 6102 45668
rect 36514 45724 36822 45733
rect 36514 45722 36520 45724
rect 36576 45722 36600 45724
rect 36656 45722 36680 45724
rect 36736 45722 36760 45724
rect 36816 45722 36822 45724
rect 36576 45670 36578 45722
rect 36758 45670 36760 45722
rect 36514 45668 36520 45670
rect 36576 45668 36600 45670
rect 36656 45668 36680 45670
rect 36736 45668 36760 45670
rect 36816 45668 36822 45670
rect 36514 45659 36822 45668
rect 67234 45724 67542 45733
rect 67234 45722 67240 45724
rect 67296 45722 67320 45724
rect 67376 45722 67400 45724
rect 67456 45722 67480 45724
rect 67536 45722 67542 45724
rect 67296 45670 67298 45722
rect 67478 45670 67480 45722
rect 67234 45668 67240 45670
rect 67296 45668 67320 45670
rect 67376 45668 67400 45670
rect 67456 45668 67480 45670
rect 67536 45668 67542 45670
rect 67234 45659 67542 45668
rect 1306 45591 1362 45600
rect 1216 41608 1268 41614
rect 1214 41576 1216 41585
rect 1268 41576 1270 41585
rect 1214 41511 1270 41520
rect 1320 38962 1348 45591
rect 5134 45180 5442 45189
rect 5134 45178 5140 45180
rect 5196 45178 5220 45180
rect 5276 45178 5300 45180
rect 5356 45178 5380 45180
rect 5436 45178 5442 45180
rect 5196 45126 5198 45178
rect 5378 45126 5380 45178
rect 5134 45124 5140 45126
rect 5196 45124 5220 45126
rect 5276 45124 5300 45126
rect 5356 45124 5380 45126
rect 5436 45124 5442 45126
rect 5134 45115 5442 45124
rect 35854 45180 36162 45189
rect 35854 45178 35860 45180
rect 35916 45178 35940 45180
rect 35996 45178 36020 45180
rect 36076 45178 36100 45180
rect 36156 45178 36162 45180
rect 35916 45126 35918 45178
rect 36098 45126 36100 45178
rect 35854 45124 35860 45126
rect 35916 45124 35940 45126
rect 35996 45124 36020 45126
rect 36076 45124 36100 45126
rect 36156 45124 36162 45126
rect 35854 45115 36162 45124
rect 66574 45180 66882 45189
rect 66574 45178 66580 45180
rect 66636 45178 66660 45180
rect 66716 45178 66740 45180
rect 66796 45178 66820 45180
rect 66876 45178 66882 45180
rect 66636 45126 66638 45178
rect 66818 45126 66820 45178
rect 66574 45124 66580 45126
rect 66636 45124 66660 45126
rect 66716 45124 66740 45126
rect 66796 45124 66820 45126
rect 66876 45124 66882 45126
rect 66574 45115 66882 45124
rect 5794 44636 6102 44645
rect 5794 44634 5800 44636
rect 5856 44634 5880 44636
rect 5936 44634 5960 44636
rect 6016 44634 6040 44636
rect 6096 44634 6102 44636
rect 5856 44582 5858 44634
rect 6038 44582 6040 44634
rect 5794 44580 5800 44582
rect 5856 44580 5880 44582
rect 5936 44580 5960 44582
rect 6016 44580 6040 44582
rect 6096 44580 6102 44582
rect 5794 44571 6102 44580
rect 36514 44636 36822 44645
rect 36514 44634 36520 44636
rect 36576 44634 36600 44636
rect 36656 44634 36680 44636
rect 36736 44634 36760 44636
rect 36816 44634 36822 44636
rect 36576 44582 36578 44634
rect 36758 44582 36760 44634
rect 36514 44580 36520 44582
rect 36576 44580 36600 44582
rect 36656 44580 36680 44582
rect 36736 44580 36760 44582
rect 36816 44580 36822 44582
rect 36514 44571 36822 44580
rect 67234 44636 67542 44645
rect 67234 44634 67240 44636
rect 67296 44634 67320 44636
rect 67376 44634 67400 44636
rect 67456 44634 67480 44636
rect 67536 44634 67542 44636
rect 67296 44582 67298 44634
rect 67478 44582 67480 44634
rect 67234 44580 67240 44582
rect 67296 44580 67320 44582
rect 67376 44580 67400 44582
rect 67456 44580 67480 44582
rect 67536 44580 67542 44582
rect 67234 44571 67542 44580
rect 5134 44092 5442 44101
rect 5134 44090 5140 44092
rect 5196 44090 5220 44092
rect 5276 44090 5300 44092
rect 5356 44090 5380 44092
rect 5436 44090 5442 44092
rect 5196 44038 5198 44090
rect 5378 44038 5380 44090
rect 5134 44036 5140 44038
rect 5196 44036 5220 44038
rect 5276 44036 5300 44038
rect 5356 44036 5380 44038
rect 5436 44036 5442 44038
rect 5134 44027 5442 44036
rect 35854 44092 36162 44101
rect 35854 44090 35860 44092
rect 35916 44090 35940 44092
rect 35996 44090 36020 44092
rect 36076 44090 36100 44092
rect 36156 44090 36162 44092
rect 35916 44038 35918 44090
rect 36098 44038 36100 44090
rect 35854 44036 35860 44038
rect 35916 44036 35940 44038
rect 35996 44036 36020 44038
rect 36076 44036 36100 44038
rect 36156 44036 36162 44038
rect 35854 44027 36162 44036
rect 66574 44092 66882 44101
rect 66574 44090 66580 44092
rect 66636 44090 66660 44092
rect 66716 44090 66740 44092
rect 66796 44090 66820 44092
rect 66876 44090 66882 44092
rect 66636 44038 66638 44090
rect 66818 44038 66820 44090
rect 66574 44036 66580 44038
rect 66636 44036 66660 44038
rect 66716 44036 66740 44038
rect 66796 44036 66820 44038
rect 66876 44036 66882 44038
rect 66574 44027 66882 44036
rect 64880 43852 64932 43858
rect 64880 43794 64932 43800
rect 5794 43548 6102 43557
rect 5794 43546 5800 43548
rect 5856 43546 5880 43548
rect 5936 43546 5960 43548
rect 6016 43546 6040 43548
rect 6096 43546 6102 43548
rect 5856 43494 5858 43546
rect 6038 43494 6040 43546
rect 5794 43492 5800 43494
rect 5856 43492 5880 43494
rect 5936 43492 5960 43494
rect 6016 43492 6040 43494
rect 6096 43492 6102 43494
rect 5794 43483 6102 43492
rect 36514 43548 36822 43557
rect 36514 43546 36520 43548
rect 36576 43546 36600 43548
rect 36656 43546 36680 43548
rect 36736 43546 36760 43548
rect 36816 43546 36822 43548
rect 36576 43494 36578 43546
rect 36758 43494 36760 43546
rect 36514 43492 36520 43494
rect 36576 43492 36600 43494
rect 36656 43492 36680 43494
rect 36736 43492 36760 43494
rect 36816 43492 36822 43494
rect 36514 43483 36822 43492
rect 5134 43004 5442 43013
rect 5134 43002 5140 43004
rect 5196 43002 5220 43004
rect 5276 43002 5300 43004
rect 5356 43002 5380 43004
rect 5436 43002 5442 43004
rect 5196 42950 5198 43002
rect 5378 42950 5380 43002
rect 5134 42948 5140 42950
rect 5196 42948 5220 42950
rect 5276 42948 5300 42950
rect 5356 42948 5380 42950
rect 5436 42948 5442 42950
rect 5134 42939 5442 42948
rect 35854 43004 36162 43013
rect 35854 43002 35860 43004
rect 35916 43002 35940 43004
rect 35996 43002 36020 43004
rect 36076 43002 36100 43004
rect 36156 43002 36162 43004
rect 35916 42950 35918 43002
rect 36098 42950 36100 43002
rect 35854 42948 35860 42950
rect 35916 42948 35940 42950
rect 35996 42948 36020 42950
rect 36076 42948 36100 42950
rect 36156 42948 36162 42950
rect 35854 42939 36162 42948
rect 60004 42764 60056 42770
rect 60004 42706 60056 42712
rect 57612 42696 57664 42702
rect 57612 42638 57664 42644
rect 5794 42460 6102 42469
rect 5794 42458 5800 42460
rect 5856 42458 5880 42460
rect 5936 42458 5960 42460
rect 6016 42458 6040 42460
rect 6096 42458 6102 42460
rect 5856 42406 5858 42458
rect 6038 42406 6040 42458
rect 5794 42404 5800 42406
rect 5856 42404 5880 42406
rect 5936 42404 5960 42406
rect 6016 42404 6040 42406
rect 6096 42404 6102 42406
rect 5794 42395 6102 42404
rect 36514 42460 36822 42469
rect 36514 42458 36520 42460
rect 36576 42458 36600 42460
rect 36656 42458 36680 42460
rect 36736 42458 36760 42460
rect 36816 42458 36822 42460
rect 36576 42406 36578 42458
rect 36758 42406 36760 42458
rect 36514 42404 36520 42406
rect 36576 42404 36600 42406
rect 36656 42404 36680 42406
rect 36736 42404 36760 42406
rect 36816 42404 36822 42406
rect 36514 42395 36822 42404
rect 5134 41916 5442 41925
rect 5134 41914 5140 41916
rect 5196 41914 5220 41916
rect 5276 41914 5300 41916
rect 5356 41914 5380 41916
rect 5436 41914 5442 41916
rect 5196 41862 5198 41914
rect 5378 41862 5380 41914
rect 5134 41860 5140 41862
rect 5196 41860 5220 41862
rect 5276 41860 5300 41862
rect 5356 41860 5380 41862
rect 5436 41860 5442 41862
rect 5134 41851 5442 41860
rect 35854 41916 36162 41925
rect 35854 41914 35860 41916
rect 35916 41914 35940 41916
rect 35996 41914 36020 41916
rect 36076 41914 36100 41916
rect 36156 41914 36162 41916
rect 35916 41862 35918 41914
rect 36098 41862 36100 41914
rect 35854 41860 35860 41862
rect 35916 41860 35940 41862
rect 35996 41860 36020 41862
rect 36076 41860 36100 41862
rect 36156 41860 36162 41862
rect 35854 41851 36162 41860
rect 5794 41372 6102 41381
rect 5794 41370 5800 41372
rect 5856 41370 5880 41372
rect 5936 41370 5960 41372
rect 6016 41370 6040 41372
rect 6096 41370 6102 41372
rect 5856 41318 5858 41370
rect 6038 41318 6040 41370
rect 5794 41316 5800 41318
rect 5856 41316 5880 41318
rect 5936 41316 5960 41318
rect 6016 41316 6040 41318
rect 6096 41316 6102 41318
rect 5794 41307 6102 41316
rect 36514 41372 36822 41381
rect 36514 41370 36520 41372
rect 36576 41370 36600 41372
rect 36656 41370 36680 41372
rect 36736 41370 36760 41372
rect 36816 41370 36822 41372
rect 36576 41318 36578 41370
rect 36758 41318 36760 41370
rect 36514 41316 36520 41318
rect 36576 41316 36600 41318
rect 36656 41316 36680 41318
rect 36736 41316 36760 41318
rect 36816 41316 36822 41318
rect 36514 41307 36822 41316
rect 5134 40828 5442 40837
rect 5134 40826 5140 40828
rect 5196 40826 5220 40828
rect 5276 40826 5300 40828
rect 5356 40826 5380 40828
rect 5436 40826 5442 40828
rect 5196 40774 5198 40826
rect 5378 40774 5380 40826
rect 5134 40772 5140 40774
rect 5196 40772 5220 40774
rect 5276 40772 5300 40774
rect 5356 40772 5380 40774
rect 5436 40772 5442 40774
rect 5134 40763 5442 40772
rect 35854 40828 36162 40837
rect 35854 40826 35860 40828
rect 35916 40826 35940 40828
rect 35996 40826 36020 40828
rect 36076 40826 36100 40828
rect 36156 40826 36162 40828
rect 35916 40774 35918 40826
rect 36098 40774 36100 40826
rect 35854 40772 35860 40774
rect 35916 40772 35940 40774
rect 35996 40772 36020 40774
rect 36076 40772 36100 40774
rect 36156 40772 36162 40774
rect 35854 40763 36162 40772
rect 57624 40458 57652 42638
rect 57980 42628 58032 42634
rect 57980 42570 58032 42576
rect 58900 42628 58952 42634
rect 58900 42570 58952 42576
rect 57992 42362 58020 42570
rect 58912 42362 58940 42570
rect 59544 42560 59596 42566
rect 59544 42502 59596 42508
rect 57980 42356 58032 42362
rect 57980 42298 58032 42304
rect 58900 42356 58952 42362
rect 58900 42298 58952 42304
rect 59556 42294 59584 42502
rect 59544 42288 59596 42294
rect 59544 42230 59596 42236
rect 58992 42220 59044 42226
rect 58992 42162 59044 42168
rect 57612 40452 57664 40458
rect 57612 40394 57664 40400
rect 5794 40284 6102 40293
rect 5794 40282 5800 40284
rect 5856 40282 5880 40284
rect 5936 40282 5960 40284
rect 6016 40282 6040 40284
rect 6096 40282 6102 40284
rect 5856 40230 5858 40282
rect 6038 40230 6040 40282
rect 5794 40228 5800 40230
rect 5856 40228 5880 40230
rect 5936 40228 5960 40230
rect 6016 40228 6040 40230
rect 6096 40228 6102 40230
rect 5794 40219 6102 40228
rect 36514 40284 36822 40293
rect 36514 40282 36520 40284
rect 36576 40282 36600 40284
rect 36656 40282 36680 40284
rect 36736 40282 36760 40284
rect 36816 40282 36822 40284
rect 36576 40230 36578 40282
rect 36758 40230 36760 40282
rect 36514 40228 36520 40230
rect 36576 40228 36600 40230
rect 36656 40228 36680 40230
rect 36736 40228 36760 40230
rect 36816 40228 36822 40230
rect 36514 40219 36822 40228
rect 5134 39740 5442 39749
rect 5134 39738 5140 39740
rect 5196 39738 5220 39740
rect 5276 39738 5300 39740
rect 5356 39738 5380 39740
rect 5436 39738 5442 39740
rect 5196 39686 5198 39738
rect 5378 39686 5380 39738
rect 5134 39684 5140 39686
rect 5196 39684 5220 39686
rect 5276 39684 5300 39686
rect 5356 39684 5380 39686
rect 5436 39684 5442 39686
rect 5134 39675 5442 39684
rect 35854 39740 36162 39749
rect 35854 39738 35860 39740
rect 35916 39738 35940 39740
rect 35996 39738 36020 39740
rect 36076 39738 36100 39740
rect 36156 39738 36162 39740
rect 35916 39686 35918 39738
rect 36098 39686 36100 39738
rect 35854 39684 35860 39686
rect 35916 39684 35940 39686
rect 35996 39684 36020 39686
rect 36076 39684 36100 39686
rect 36156 39684 36162 39686
rect 35854 39675 36162 39684
rect 57624 39506 57652 40394
rect 59004 40050 59032 42162
rect 58992 40044 59044 40050
rect 58992 39986 59044 39992
rect 57612 39500 57664 39506
rect 57612 39442 57664 39448
rect 59004 39438 59032 39986
rect 58348 39432 58400 39438
rect 58348 39374 58400 39380
rect 58992 39432 59044 39438
rect 58992 39374 59044 39380
rect 57060 39364 57112 39370
rect 57060 39306 57112 39312
rect 5794 39196 6102 39205
rect 5794 39194 5800 39196
rect 5856 39194 5880 39196
rect 5936 39194 5960 39196
rect 6016 39194 6040 39196
rect 6096 39194 6102 39196
rect 5856 39142 5858 39194
rect 6038 39142 6040 39194
rect 5794 39140 5800 39142
rect 5856 39140 5880 39142
rect 5936 39140 5960 39142
rect 6016 39140 6040 39142
rect 6096 39140 6102 39142
rect 5794 39131 6102 39140
rect 36514 39196 36822 39205
rect 36514 39194 36520 39196
rect 36576 39194 36600 39196
rect 36656 39194 36680 39196
rect 36736 39194 36760 39196
rect 36816 39194 36822 39196
rect 36576 39142 36578 39194
rect 36758 39142 36760 39194
rect 36514 39140 36520 39142
rect 36576 39140 36600 39142
rect 36656 39140 36680 39142
rect 36736 39140 36760 39142
rect 36816 39140 36822 39142
rect 36514 39131 36822 39140
rect 1308 38956 1360 38962
rect 1308 38898 1360 38904
rect 5134 38652 5442 38661
rect 5134 38650 5140 38652
rect 5196 38650 5220 38652
rect 5276 38650 5300 38652
rect 5356 38650 5380 38652
rect 5436 38650 5442 38652
rect 5196 38598 5198 38650
rect 5378 38598 5380 38650
rect 5134 38596 5140 38598
rect 5196 38596 5220 38598
rect 5276 38596 5300 38598
rect 5356 38596 5380 38598
rect 5436 38596 5442 38598
rect 5134 38587 5442 38596
rect 35854 38652 36162 38661
rect 35854 38650 35860 38652
rect 35916 38650 35940 38652
rect 35996 38650 36020 38652
rect 36076 38650 36100 38652
rect 36156 38650 36162 38652
rect 35916 38598 35918 38650
rect 36098 38598 36100 38650
rect 35854 38596 35860 38598
rect 35916 38596 35940 38598
rect 35996 38596 36020 38598
rect 36076 38596 36100 38598
rect 36156 38596 36162 38598
rect 35854 38587 36162 38596
rect 57072 38554 57100 39306
rect 57980 39296 58032 39302
rect 57980 39238 58032 39244
rect 57060 38548 57112 38554
rect 57060 38490 57112 38496
rect 57336 38344 57388 38350
rect 57336 38286 57388 38292
rect 5794 38108 6102 38117
rect 5794 38106 5800 38108
rect 5856 38106 5880 38108
rect 5936 38106 5960 38108
rect 6016 38106 6040 38108
rect 6096 38106 6102 38108
rect 5856 38054 5858 38106
rect 6038 38054 6040 38106
rect 5794 38052 5800 38054
rect 5856 38052 5880 38054
rect 5936 38052 5960 38054
rect 6016 38052 6040 38054
rect 6096 38052 6102 38054
rect 5794 38043 6102 38052
rect 36514 38108 36822 38117
rect 36514 38106 36520 38108
rect 36576 38106 36600 38108
rect 36656 38106 36680 38108
rect 36736 38106 36760 38108
rect 36816 38106 36822 38108
rect 36576 38054 36578 38106
rect 36758 38054 36760 38106
rect 36514 38052 36520 38054
rect 36576 38052 36600 38054
rect 36656 38052 36680 38054
rect 36736 38052 36760 38054
rect 36816 38052 36822 38054
rect 36514 38043 36822 38052
rect 5134 37564 5442 37573
rect 5134 37562 5140 37564
rect 5196 37562 5220 37564
rect 5276 37562 5300 37564
rect 5356 37562 5380 37564
rect 5436 37562 5442 37564
rect 5196 37510 5198 37562
rect 5378 37510 5380 37562
rect 5134 37508 5140 37510
rect 5196 37508 5220 37510
rect 5276 37508 5300 37510
rect 5356 37508 5380 37510
rect 5436 37508 5442 37510
rect 5134 37499 5442 37508
rect 35854 37564 36162 37573
rect 35854 37562 35860 37564
rect 35916 37562 35940 37564
rect 35996 37562 36020 37564
rect 36076 37562 36100 37564
rect 36156 37562 36162 37564
rect 35916 37510 35918 37562
rect 36098 37510 36100 37562
rect 35854 37508 35860 37510
rect 35916 37508 35940 37510
rect 35996 37508 36020 37510
rect 36076 37508 36100 37510
rect 36156 37508 36162 37510
rect 35854 37499 36162 37508
rect 57348 37126 57376 38286
rect 57992 38282 58020 39238
rect 57796 38276 57848 38282
rect 57796 38218 57848 38224
rect 57980 38276 58032 38282
rect 57980 38218 58032 38224
rect 57808 37262 57836 38218
rect 57796 37256 57848 37262
rect 57796 37198 57848 37204
rect 57992 37194 58020 38218
rect 57980 37188 58032 37194
rect 57980 37130 58032 37136
rect 56784 37120 56836 37126
rect 56784 37062 56836 37068
rect 57336 37120 57388 37126
rect 57336 37062 57388 37068
rect 5794 37020 6102 37029
rect 5794 37018 5800 37020
rect 5856 37018 5880 37020
rect 5936 37018 5960 37020
rect 6016 37018 6040 37020
rect 6096 37018 6102 37020
rect 5856 36966 5858 37018
rect 6038 36966 6040 37018
rect 5794 36964 5800 36966
rect 5856 36964 5880 36966
rect 5936 36964 5960 36966
rect 6016 36964 6040 36966
rect 6096 36964 6102 36966
rect 5794 36955 6102 36964
rect 36514 37020 36822 37029
rect 36514 37018 36520 37020
rect 36576 37018 36600 37020
rect 36656 37018 36680 37020
rect 36736 37018 36760 37020
rect 36816 37018 36822 37020
rect 36576 36966 36578 37018
rect 36758 36966 36760 37018
rect 36514 36964 36520 36966
rect 36576 36964 36600 36966
rect 36656 36964 36680 36966
rect 36736 36964 36760 36966
rect 36816 36964 36822 36966
rect 36514 36955 36822 36964
rect 5134 36476 5442 36485
rect 5134 36474 5140 36476
rect 5196 36474 5220 36476
rect 5276 36474 5300 36476
rect 5356 36474 5380 36476
rect 5436 36474 5442 36476
rect 5196 36422 5198 36474
rect 5378 36422 5380 36474
rect 5134 36420 5140 36422
rect 5196 36420 5220 36422
rect 5276 36420 5300 36422
rect 5356 36420 5380 36422
rect 5436 36420 5442 36422
rect 5134 36411 5442 36420
rect 35854 36476 36162 36485
rect 35854 36474 35860 36476
rect 35916 36474 35940 36476
rect 35996 36474 36020 36476
rect 36076 36474 36100 36476
rect 36156 36474 36162 36476
rect 35916 36422 35918 36474
rect 36098 36422 36100 36474
rect 35854 36420 35860 36422
rect 35916 36420 35940 36422
rect 35996 36420 36020 36422
rect 36076 36420 36100 36422
rect 36156 36420 36162 36422
rect 35854 36411 36162 36420
rect 5794 35932 6102 35941
rect 5794 35930 5800 35932
rect 5856 35930 5880 35932
rect 5936 35930 5960 35932
rect 6016 35930 6040 35932
rect 6096 35930 6102 35932
rect 5856 35878 5858 35930
rect 6038 35878 6040 35930
rect 5794 35876 5800 35878
rect 5856 35876 5880 35878
rect 5936 35876 5960 35878
rect 6016 35876 6040 35878
rect 6096 35876 6102 35878
rect 5794 35867 6102 35876
rect 36514 35932 36822 35941
rect 36514 35930 36520 35932
rect 36576 35930 36600 35932
rect 36656 35930 36680 35932
rect 36736 35930 36760 35932
rect 36816 35930 36822 35932
rect 36576 35878 36578 35930
rect 36758 35878 36760 35930
rect 36514 35876 36520 35878
rect 36576 35876 36600 35878
rect 36656 35876 36680 35878
rect 36736 35876 36760 35878
rect 36816 35876 36822 35878
rect 36514 35867 36822 35876
rect 56796 35630 56824 37062
rect 57992 36786 58020 37130
rect 57980 36780 58032 36786
rect 57980 36722 58032 36728
rect 58072 35692 58124 35698
rect 58072 35634 58124 35640
rect 56784 35624 56836 35630
rect 56784 35566 56836 35572
rect 1216 35488 1268 35494
rect 1214 35456 1216 35465
rect 56416 35488 56468 35494
rect 1268 35456 1270 35465
rect 56416 35430 56468 35436
rect 1214 35391 1270 35400
rect 5134 35388 5442 35397
rect 5134 35386 5140 35388
rect 5196 35386 5220 35388
rect 5276 35386 5300 35388
rect 5356 35386 5380 35388
rect 5436 35386 5442 35388
rect 5196 35334 5198 35386
rect 5378 35334 5380 35386
rect 5134 35332 5140 35334
rect 5196 35332 5220 35334
rect 5276 35332 5300 35334
rect 5356 35332 5380 35334
rect 5436 35332 5442 35334
rect 5134 35323 5442 35332
rect 35854 35388 36162 35397
rect 35854 35386 35860 35388
rect 35916 35386 35940 35388
rect 35996 35386 36020 35388
rect 36076 35386 36100 35388
rect 36156 35386 36162 35388
rect 35916 35334 35918 35386
rect 36098 35334 36100 35386
rect 35854 35332 35860 35334
rect 35916 35332 35940 35334
rect 35996 35332 36020 35334
rect 36076 35332 36100 35334
rect 36156 35332 36162 35334
rect 35854 35323 36162 35332
rect 56428 35290 56456 35430
rect 58084 35290 58112 35634
rect 58360 35562 58388 39374
rect 60016 37262 60044 42706
rect 64892 41818 64920 43794
rect 66904 43784 66956 43790
rect 66904 43726 66956 43732
rect 65432 43648 65484 43654
rect 65432 43590 65484 43596
rect 65444 43382 65472 43590
rect 66916 43450 66944 43726
rect 67234 43548 67542 43557
rect 67234 43546 67240 43548
rect 67296 43546 67320 43548
rect 67376 43546 67400 43548
rect 67456 43546 67480 43548
rect 67536 43546 67542 43548
rect 67296 43494 67298 43546
rect 67478 43494 67480 43546
rect 67234 43492 67240 43494
rect 67296 43492 67320 43494
rect 67376 43492 67400 43494
rect 67456 43492 67480 43494
rect 67536 43492 67542 43494
rect 67234 43483 67542 43492
rect 66260 43444 66312 43450
rect 66260 43386 66312 43392
rect 66904 43444 66956 43450
rect 66904 43386 66956 43392
rect 65432 43376 65484 43382
rect 65432 43318 65484 43324
rect 65156 43240 65208 43246
rect 65156 43182 65208 43188
rect 64880 41812 64932 41818
rect 64880 41754 64932 41760
rect 64604 41608 64656 41614
rect 64604 41550 64656 41556
rect 64788 41608 64840 41614
rect 64788 41550 64840 41556
rect 62672 40656 62724 40662
rect 62672 40598 62724 40604
rect 60924 40588 60976 40594
rect 60924 40530 60976 40536
rect 60832 40520 60884 40526
rect 60832 40462 60884 40468
rect 60844 40186 60872 40462
rect 60936 40390 60964 40530
rect 62120 40452 62172 40458
rect 62120 40394 62172 40400
rect 60924 40384 60976 40390
rect 60924 40326 60976 40332
rect 60832 40180 60884 40186
rect 60832 40122 60884 40128
rect 60004 37256 60056 37262
rect 60004 37198 60056 37204
rect 60016 36854 60044 37198
rect 60936 36854 60964 40326
rect 62132 40050 62160 40394
rect 62684 40050 62712 40598
rect 63500 40588 63552 40594
rect 63500 40530 63552 40536
rect 62120 40044 62172 40050
rect 62120 39986 62172 39992
rect 62672 40044 62724 40050
rect 62672 39986 62724 39992
rect 63512 38554 63540 40530
rect 64616 40390 64644 41550
rect 64800 40662 64828 41550
rect 64788 40656 64840 40662
rect 64788 40598 64840 40604
rect 64800 40526 64828 40598
rect 65168 40594 65196 43182
rect 66272 40746 66300 43386
rect 67088 43240 67140 43246
rect 67088 43182 67140 43188
rect 66574 43004 66882 43013
rect 66574 43002 66580 43004
rect 66636 43002 66660 43004
rect 66716 43002 66740 43004
rect 66796 43002 66820 43004
rect 66876 43002 66882 43004
rect 66636 42950 66638 43002
rect 66818 42950 66820 43002
rect 66574 42948 66580 42950
rect 66636 42948 66660 42950
rect 66716 42948 66740 42950
rect 66796 42948 66820 42950
rect 66876 42948 66882 42950
rect 66574 42939 66882 42948
rect 66574 41916 66882 41925
rect 66574 41914 66580 41916
rect 66636 41914 66660 41916
rect 66716 41914 66740 41916
rect 66796 41914 66820 41916
rect 66876 41914 66882 41916
rect 66636 41862 66638 41914
rect 66818 41862 66820 41914
rect 66574 41860 66580 41862
rect 66636 41860 66660 41862
rect 66716 41860 66740 41862
rect 66796 41860 66820 41862
rect 66876 41860 66882 41862
rect 66574 41851 66882 41860
rect 66574 40828 66882 40837
rect 66574 40826 66580 40828
rect 66636 40826 66660 40828
rect 66716 40826 66740 40828
rect 66796 40826 66820 40828
rect 66876 40826 66882 40828
rect 66636 40774 66638 40826
rect 66818 40774 66820 40826
rect 66574 40772 66580 40774
rect 66636 40772 66660 40774
rect 66716 40772 66740 40774
rect 66796 40772 66820 40774
rect 66876 40772 66882 40774
rect 66574 40763 66882 40772
rect 66088 40718 66300 40746
rect 66088 40610 66116 40718
rect 65156 40588 65208 40594
rect 65156 40530 65208 40536
rect 65996 40582 66116 40610
rect 66168 40588 66220 40594
rect 65996 40526 66024 40582
rect 66168 40530 66220 40536
rect 64788 40520 64840 40526
rect 64788 40462 64840 40468
rect 65984 40520 66036 40526
rect 65984 40462 66036 40468
rect 66076 40520 66128 40526
rect 66076 40462 66128 40468
rect 64604 40384 64656 40390
rect 64604 40326 64656 40332
rect 64616 40186 64644 40326
rect 64604 40180 64656 40186
rect 64604 40122 64656 40128
rect 65996 40050 66024 40462
rect 66088 40186 66116 40462
rect 66076 40180 66128 40186
rect 66076 40122 66128 40128
rect 66180 40118 66208 40530
rect 66168 40112 66220 40118
rect 66168 40054 66220 40060
rect 65984 40044 66036 40050
rect 65984 39986 66036 39992
rect 65800 39840 65852 39846
rect 65800 39782 65852 39788
rect 63500 38548 63552 38554
rect 63500 38490 63552 38496
rect 63512 37330 63540 38490
rect 63500 37324 63552 37330
rect 63500 37266 63552 37272
rect 65340 37324 65392 37330
rect 65340 37266 65392 37272
rect 60004 36848 60056 36854
rect 60004 36790 60056 36796
rect 60372 36848 60424 36854
rect 60372 36790 60424 36796
rect 60924 36848 60976 36854
rect 60924 36790 60976 36796
rect 60016 36310 60044 36790
rect 60188 36780 60240 36786
rect 60188 36722 60240 36728
rect 60280 36780 60332 36786
rect 60280 36722 60332 36728
rect 60004 36304 60056 36310
rect 60004 36246 60056 36252
rect 60200 36242 60228 36722
rect 60292 36242 60320 36722
rect 60188 36236 60240 36242
rect 60188 36178 60240 36184
rect 60280 36236 60332 36242
rect 60280 36178 60332 36184
rect 60292 35698 60320 36178
rect 60384 36106 60412 36790
rect 60936 36242 60964 36790
rect 60924 36236 60976 36242
rect 60924 36178 60976 36184
rect 60372 36100 60424 36106
rect 60372 36042 60424 36048
rect 60556 36032 60608 36038
rect 60556 35974 60608 35980
rect 62120 36032 62172 36038
rect 62120 35974 62172 35980
rect 60568 35766 60596 35974
rect 60556 35760 60608 35766
rect 60556 35702 60608 35708
rect 60280 35692 60332 35698
rect 60280 35634 60332 35640
rect 62132 35630 62160 35974
rect 63512 35834 63540 37266
rect 65352 36922 65380 37266
rect 65340 36916 65392 36922
rect 65340 36858 65392 36864
rect 65812 36786 65840 39782
rect 66180 39574 66208 40054
rect 66168 39568 66220 39574
rect 66168 39510 66220 39516
rect 66272 39438 66300 40718
rect 66904 40656 66956 40662
rect 66904 40598 66956 40604
rect 66444 40384 66496 40390
rect 66444 40326 66496 40332
rect 66456 39914 66484 40326
rect 66916 40050 66944 40598
rect 66996 40452 67048 40458
rect 66996 40394 67048 40400
rect 67008 40050 67036 40394
rect 66904 40044 66956 40050
rect 66904 39986 66956 39992
rect 66996 40044 67048 40050
rect 66996 39986 67048 39992
rect 66444 39908 66496 39914
rect 66444 39850 66496 39856
rect 66574 39740 66882 39749
rect 66574 39738 66580 39740
rect 66636 39738 66660 39740
rect 66716 39738 66740 39740
rect 66796 39738 66820 39740
rect 66876 39738 66882 39740
rect 66636 39686 66638 39738
rect 66818 39686 66820 39738
rect 66574 39684 66580 39686
rect 66636 39684 66660 39686
rect 66716 39684 66740 39686
rect 66796 39684 66820 39686
rect 66876 39684 66882 39686
rect 66574 39675 66882 39684
rect 66916 39438 66944 39986
rect 67100 39982 67128 43182
rect 67234 42460 67542 42469
rect 67234 42458 67240 42460
rect 67296 42458 67320 42460
rect 67376 42458 67400 42460
rect 67456 42458 67480 42460
rect 67536 42458 67542 42460
rect 67296 42406 67298 42458
rect 67478 42406 67480 42458
rect 67234 42404 67240 42406
rect 67296 42404 67320 42406
rect 67376 42404 67400 42406
rect 67456 42404 67480 42406
rect 67536 42404 67542 42406
rect 67234 42395 67542 42404
rect 74356 41608 74408 41614
rect 74356 41550 74408 41556
rect 76380 41608 76432 41614
rect 76380 41550 76432 41556
rect 71228 41472 71280 41478
rect 71228 41414 71280 41420
rect 67234 41372 67542 41381
rect 67234 41370 67240 41372
rect 67296 41370 67320 41372
rect 67376 41370 67400 41372
rect 67456 41370 67480 41372
rect 67536 41370 67542 41372
rect 67296 41318 67298 41370
rect 67478 41318 67480 41370
rect 67234 41316 67240 41318
rect 67296 41316 67320 41318
rect 67376 41316 67400 41318
rect 67456 41316 67480 41318
rect 67536 41316 67542 41318
rect 67234 41307 67542 41316
rect 71240 41206 71268 41414
rect 74368 41274 74396 41550
rect 74632 41540 74684 41546
rect 74632 41482 74684 41488
rect 74356 41268 74408 41274
rect 74356 41210 74408 41216
rect 71228 41200 71280 41206
rect 71228 41142 71280 41148
rect 68284 41132 68336 41138
rect 68284 41074 68336 41080
rect 68296 40594 68324 41074
rect 74644 41070 74672 41482
rect 75920 41472 75972 41478
rect 75920 41414 75972 41420
rect 75932 41070 75960 41414
rect 70492 41064 70544 41070
rect 70492 41006 70544 41012
rect 71136 41064 71188 41070
rect 71136 41006 71188 41012
rect 74632 41064 74684 41070
rect 74632 41006 74684 41012
rect 75920 41064 75972 41070
rect 75920 41006 75972 41012
rect 70504 40730 70532 41006
rect 70492 40724 70544 40730
rect 70492 40666 70544 40672
rect 71148 40594 71176 41006
rect 71964 40928 72016 40934
rect 71964 40870 72016 40876
rect 71504 40656 71556 40662
rect 71504 40598 71556 40604
rect 68284 40588 68336 40594
rect 68284 40530 68336 40536
rect 71136 40588 71188 40594
rect 71136 40530 71188 40536
rect 68008 40452 68060 40458
rect 68008 40394 68060 40400
rect 67234 40284 67542 40293
rect 67234 40282 67240 40284
rect 67296 40282 67320 40284
rect 67376 40282 67400 40284
rect 67456 40282 67480 40284
rect 67536 40282 67542 40284
rect 67296 40230 67298 40282
rect 67478 40230 67480 40282
rect 67234 40228 67240 40230
rect 67296 40228 67320 40230
rect 67376 40228 67400 40230
rect 67456 40228 67480 40230
rect 67536 40228 67542 40230
rect 67234 40219 67542 40228
rect 68020 40186 68048 40394
rect 68008 40180 68060 40186
rect 68008 40122 68060 40128
rect 67088 39976 67140 39982
rect 67088 39918 67140 39924
rect 66260 39432 66312 39438
rect 66260 39374 66312 39380
rect 66904 39432 66956 39438
rect 67100 39386 67128 39918
rect 66904 39374 66956 39380
rect 67008 39358 67128 39386
rect 66904 39296 66956 39302
rect 66904 39238 66956 39244
rect 66444 38752 66496 38758
rect 66444 38694 66496 38700
rect 66456 38282 66484 38694
rect 66574 38652 66882 38661
rect 66574 38650 66580 38652
rect 66636 38650 66660 38652
rect 66716 38650 66740 38652
rect 66796 38650 66820 38652
rect 66876 38650 66882 38652
rect 66636 38598 66638 38650
rect 66818 38598 66820 38650
rect 66574 38596 66580 38598
rect 66636 38596 66660 38598
rect 66716 38596 66740 38598
rect 66796 38596 66820 38598
rect 66876 38596 66882 38598
rect 66574 38587 66882 38596
rect 66444 38276 66496 38282
rect 66444 38218 66496 38224
rect 66574 37564 66882 37573
rect 66574 37562 66580 37564
rect 66636 37562 66660 37564
rect 66716 37562 66740 37564
rect 66796 37562 66820 37564
rect 66876 37562 66882 37564
rect 66636 37510 66638 37562
rect 66818 37510 66820 37562
rect 66574 37508 66580 37510
rect 66636 37508 66660 37510
rect 66716 37508 66740 37510
rect 66796 37508 66820 37510
rect 66876 37508 66882 37510
rect 66574 37499 66882 37508
rect 66916 37262 66944 39238
rect 66904 37256 66956 37262
rect 66904 37198 66956 37204
rect 65984 37188 66036 37194
rect 65984 37130 66036 37136
rect 65996 36922 66024 37130
rect 66536 37120 66588 37126
rect 66536 37062 66588 37068
rect 65984 36916 66036 36922
rect 65984 36858 66036 36864
rect 66548 36854 66576 37062
rect 66536 36848 66588 36854
rect 66536 36790 66588 36796
rect 67008 36786 67036 39358
rect 67088 39296 67140 39302
rect 67088 39238 67140 39244
rect 65616 36780 65668 36786
rect 65616 36722 65668 36728
rect 65800 36780 65852 36786
rect 65800 36722 65852 36728
rect 66168 36780 66220 36786
rect 66168 36722 66220 36728
rect 66996 36780 67048 36786
rect 66996 36722 67048 36728
rect 65628 36378 65656 36722
rect 65616 36372 65668 36378
rect 65616 36314 65668 36320
rect 65984 36372 66036 36378
rect 65984 36314 66036 36320
rect 63500 35828 63552 35834
rect 63500 35770 63552 35776
rect 60372 35624 60424 35630
rect 60372 35566 60424 35572
rect 62120 35624 62172 35630
rect 62120 35566 62172 35572
rect 58348 35556 58400 35562
rect 58348 35498 58400 35504
rect 56416 35284 56468 35290
rect 56416 35226 56468 35232
rect 58072 35284 58124 35290
rect 58072 35226 58124 35232
rect 58360 35086 58388 35498
rect 60384 35154 60412 35566
rect 60372 35148 60424 35154
rect 60372 35090 60424 35096
rect 58348 35080 58400 35086
rect 58348 35022 58400 35028
rect 5794 34844 6102 34853
rect 5794 34842 5800 34844
rect 5856 34842 5880 34844
rect 5936 34842 5960 34844
rect 6016 34842 6040 34844
rect 6096 34842 6102 34844
rect 5856 34790 5858 34842
rect 6038 34790 6040 34842
rect 5794 34788 5800 34790
rect 5856 34788 5880 34790
rect 5936 34788 5960 34790
rect 6016 34788 6040 34790
rect 6096 34788 6102 34790
rect 5794 34779 6102 34788
rect 36514 34844 36822 34853
rect 36514 34842 36520 34844
rect 36576 34842 36600 34844
rect 36656 34842 36680 34844
rect 36736 34842 36760 34844
rect 36816 34842 36822 34844
rect 36576 34790 36578 34842
rect 36758 34790 36760 34842
rect 36514 34788 36520 34790
rect 36576 34788 36600 34790
rect 36656 34788 36680 34790
rect 36736 34788 36760 34790
rect 36816 34788 36822 34790
rect 36514 34779 36822 34788
rect 65996 34542 66024 36314
rect 66180 35698 66208 36722
rect 66574 36476 66882 36485
rect 66574 36474 66580 36476
rect 66636 36474 66660 36476
rect 66716 36474 66740 36476
rect 66796 36474 66820 36476
rect 66876 36474 66882 36476
rect 66636 36422 66638 36474
rect 66818 36422 66820 36474
rect 66574 36420 66580 36422
rect 66636 36420 66660 36422
rect 66716 36420 66740 36422
rect 66796 36420 66820 36422
rect 66876 36420 66882 36422
rect 66574 36411 66882 36420
rect 67100 36174 67128 39238
rect 67234 39196 67542 39205
rect 67234 39194 67240 39196
rect 67296 39194 67320 39196
rect 67376 39194 67400 39196
rect 67456 39194 67480 39196
rect 67536 39194 67542 39196
rect 67296 39142 67298 39194
rect 67478 39142 67480 39194
rect 67234 39140 67240 39142
rect 67296 39140 67320 39142
rect 67376 39140 67400 39142
rect 67456 39140 67480 39142
rect 67536 39140 67542 39142
rect 67234 39131 67542 39140
rect 68296 38554 68324 40530
rect 71148 39642 71176 40530
rect 71136 39636 71188 39642
rect 71136 39578 71188 39584
rect 70676 39364 70728 39370
rect 70676 39306 70728 39312
rect 70688 38894 70716 39306
rect 71044 39296 71096 39302
rect 71044 39238 71096 39244
rect 71228 39296 71280 39302
rect 71228 39238 71280 39244
rect 71056 38962 71084 39238
rect 71240 39114 71268 39238
rect 71148 39098 71268 39114
rect 71516 39098 71544 40598
rect 71596 39364 71648 39370
rect 71596 39306 71648 39312
rect 71608 39098 71636 39306
rect 71136 39092 71268 39098
rect 71188 39086 71268 39092
rect 71504 39092 71556 39098
rect 71136 39034 71188 39040
rect 71504 39034 71556 39040
rect 71596 39092 71648 39098
rect 71596 39034 71648 39040
rect 71044 38956 71096 38962
rect 71044 38898 71096 38904
rect 70676 38888 70728 38894
rect 70676 38830 70728 38836
rect 68284 38548 68336 38554
rect 68284 38490 68336 38496
rect 68928 38548 68980 38554
rect 68928 38490 68980 38496
rect 67234 38108 67542 38117
rect 67234 38106 67240 38108
rect 67296 38106 67320 38108
rect 67376 38106 67400 38108
rect 67456 38106 67480 38108
rect 67536 38106 67542 38108
rect 67296 38054 67298 38106
rect 67478 38054 67480 38106
rect 67234 38052 67240 38054
rect 67296 38052 67320 38054
rect 67376 38052 67400 38054
rect 67456 38052 67480 38054
rect 67536 38052 67542 38054
rect 67234 38043 67542 38052
rect 68296 37942 68324 38490
rect 68284 37936 68336 37942
rect 68284 37878 68336 37884
rect 67234 37020 67542 37029
rect 67234 37018 67240 37020
rect 67296 37018 67320 37020
rect 67376 37018 67400 37020
rect 67456 37018 67480 37020
rect 67536 37018 67542 37020
rect 67296 36966 67298 37018
rect 67478 36966 67480 37018
rect 67234 36964 67240 36966
rect 67296 36964 67320 36966
rect 67376 36964 67400 36966
rect 67456 36964 67480 36966
rect 67536 36964 67542 36966
rect 67234 36955 67542 36964
rect 67088 36168 67140 36174
rect 67088 36110 67140 36116
rect 67234 35932 67542 35941
rect 67234 35930 67240 35932
rect 67296 35930 67320 35932
rect 67376 35930 67400 35932
rect 67456 35930 67480 35932
rect 67536 35930 67542 35932
rect 67296 35878 67298 35930
rect 67478 35878 67480 35930
rect 67234 35876 67240 35878
rect 67296 35876 67320 35878
rect 67376 35876 67400 35878
rect 67456 35876 67480 35878
rect 67536 35876 67542 35878
rect 67234 35867 67542 35876
rect 66168 35692 66220 35698
rect 66168 35634 66220 35640
rect 66180 34626 66208 35634
rect 66574 35388 66882 35397
rect 66574 35386 66580 35388
rect 66636 35386 66660 35388
rect 66716 35386 66740 35388
rect 66796 35386 66820 35388
rect 66876 35386 66882 35388
rect 66636 35334 66638 35386
rect 66818 35334 66820 35386
rect 66574 35332 66580 35334
rect 66636 35332 66660 35334
rect 66716 35332 66740 35334
rect 66796 35332 66820 35334
rect 66876 35332 66882 35334
rect 66574 35323 66882 35332
rect 66996 35080 67048 35086
rect 66996 35022 67048 35028
rect 66180 34598 66300 34626
rect 67008 34610 67036 35022
rect 67234 34844 67542 34853
rect 67234 34842 67240 34844
rect 67296 34842 67320 34844
rect 67376 34842 67400 34844
rect 67456 34842 67480 34844
rect 67536 34842 67542 34844
rect 67296 34790 67298 34842
rect 67478 34790 67480 34842
rect 67234 34788 67240 34790
rect 67296 34788 67320 34790
rect 67376 34788 67400 34790
rect 67456 34788 67480 34790
rect 67536 34788 67542 34790
rect 67234 34779 67542 34788
rect 68940 34746 68968 38490
rect 70688 36106 70716 38830
rect 71056 36174 71084 38898
rect 70860 36168 70912 36174
rect 70860 36110 70912 36116
rect 71044 36168 71096 36174
rect 71044 36110 71096 36116
rect 70676 36100 70728 36106
rect 70676 36042 70728 36048
rect 70688 35766 70716 36042
rect 70676 35760 70728 35766
rect 70676 35702 70728 35708
rect 70124 35624 70176 35630
rect 70124 35566 70176 35572
rect 70136 35154 70164 35566
rect 70676 35556 70728 35562
rect 70676 35498 70728 35504
rect 70124 35148 70176 35154
rect 70124 35090 70176 35096
rect 68928 34740 68980 34746
rect 68928 34682 68980 34688
rect 65984 34536 66036 34542
rect 65984 34478 66036 34484
rect 5134 34300 5442 34309
rect 5134 34298 5140 34300
rect 5196 34298 5220 34300
rect 5276 34298 5300 34300
rect 5356 34298 5380 34300
rect 5436 34298 5442 34300
rect 5196 34246 5198 34298
rect 5378 34246 5380 34298
rect 5134 34244 5140 34246
rect 5196 34244 5220 34246
rect 5276 34244 5300 34246
rect 5356 34244 5380 34246
rect 5436 34244 5442 34246
rect 5134 34235 5442 34244
rect 35854 34300 36162 34309
rect 35854 34298 35860 34300
rect 35916 34298 35940 34300
rect 35996 34298 36020 34300
rect 36076 34298 36100 34300
rect 36156 34298 36162 34300
rect 35916 34246 35918 34298
rect 36098 34246 36100 34298
rect 35854 34244 35860 34246
rect 35916 34244 35940 34246
rect 35996 34244 36020 34246
rect 36076 34244 36100 34246
rect 36156 34244 36162 34246
rect 35854 34235 36162 34244
rect 66272 33862 66300 34598
rect 66996 34604 67048 34610
rect 66996 34546 67048 34552
rect 66574 34300 66882 34309
rect 66574 34298 66580 34300
rect 66636 34298 66660 34300
rect 66716 34298 66740 34300
rect 66796 34298 66820 34300
rect 66876 34298 66882 34300
rect 66636 34246 66638 34298
rect 66818 34246 66820 34298
rect 66574 34244 66580 34246
rect 66636 34244 66660 34246
rect 66716 34244 66740 34246
rect 66796 34244 66820 34246
rect 66876 34244 66882 34246
rect 66574 34235 66882 34244
rect 67008 34202 67036 34546
rect 68008 34400 68060 34406
rect 68008 34342 68060 34348
rect 66996 34196 67048 34202
rect 66996 34138 67048 34144
rect 68020 34066 68048 34342
rect 68940 34066 68968 34682
rect 70136 34542 70164 35090
rect 70688 35086 70716 35498
rect 70872 35290 70900 36110
rect 71148 36106 71176 39034
rect 71976 38962 72004 40870
rect 75736 39432 75788 39438
rect 75736 39374 75788 39380
rect 71964 38956 72016 38962
rect 71964 38898 72016 38904
rect 74632 38956 74684 38962
rect 74632 38898 74684 38904
rect 74644 38350 74672 38898
rect 75748 38894 75776 39374
rect 75828 39364 75880 39370
rect 75828 39306 75880 39312
rect 75736 38888 75788 38894
rect 75736 38830 75788 38836
rect 75368 38752 75420 38758
rect 75368 38694 75420 38700
rect 74632 38344 74684 38350
rect 74632 38286 74684 38292
rect 75380 37262 75408 38694
rect 75748 38570 75776 38830
rect 75840 38758 75868 39306
rect 75932 39098 75960 41006
rect 76196 39568 76248 39574
rect 76196 39510 76248 39516
rect 76012 39296 76064 39302
rect 76012 39238 76064 39244
rect 75920 39092 75972 39098
rect 75920 39034 75972 39040
rect 75828 38752 75880 38758
rect 75828 38694 75880 38700
rect 75748 38542 75868 38570
rect 76024 38554 76052 39238
rect 75368 37256 75420 37262
rect 75368 37198 75420 37204
rect 71688 36236 71740 36242
rect 71688 36178 71740 36184
rect 71136 36100 71188 36106
rect 71136 36042 71188 36048
rect 71148 35698 71176 36042
rect 71700 35698 71728 36178
rect 73160 36168 73212 36174
rect 73160 36110 73212 36116
rect 74080 36168 74132 36174
rect 74080 36110 74132 36116
rect 73172 35834 73200 36110
rect 73160 35828 73212 35834
rect 73160 35770 73212 35776
rect 71136 35692 71188 35698
rect 71136 35634 71188 35640
rect 71688 35692 71740 35698
rect 71688 35634 71740 35640
rect 71320 35488 71372 35494
rect 71320 35430 71372 35436
rect 70860 35284 70912 35290
rect 70860 35226 70912 35232
rect 70676 35080 70728 35086
rect 70676 35022 70728 35028
rect 71332 34678 71360 35430
rect 74092 34678 74120 36110
rect 75840 36038 75868 38542
rect 76012 38548 76064 38554
rect 76012 38490 76064 38496
rect 76208 38434 76236 39510
rect 76288 38956 76340 38962
rect 76288 38898 76340 38904
rect 76300 38554 76328 38898
rect 76288 38548 76340 38554
rect 76288 38490 76340 38496
rect 76208 38406 76328 38434
rect 76300 38350 76328 38406
rect 76104 38344 76156 38350
rect 76104 38286 76156 38292
rect 76288 38344 76340 38350
rect 76288 38286 76340 38292
rect 76116 37194 76144 38286
rect 76104 37188 76156 37194
rect 76104 37130 76156 37136
rect 76300 36174 76328 38286
rect 76392 36242 76420 41550
rect 77482 38856 77538 38865
rect 77482 38791 77484 38800
rect 77536 38791 77538 38800
rect 77484 38762 77536 38768
rect 77484 38208 77536 38214
rect 77482 38176 77484 38185
rect 77536 38176 77538 38185
rect 77482 38111 77538 38120
rect 76472 37868 76524 37874
rect 76472 37810 76524 37816
rect 76484 36378 76512 37810
rect 77484 37664 77536 37670
rect 77484 37606 77536 37612
rect 77496 37505 77524 37606
rect 77482 37496 77538 37505
rect 77482 37431 77538 37440
rect 77484 37120 77536 37126
rect 77484 37062 77536 37068
rect 77496 36825 77524 37062
rect 77482 36816 77538 36825
rect 77482 36751 77538 36760
rect 76472 36372 76524 36378
rect 76472 36314 76524 36320
rect 76380 36236 76432 36242
rect 76380 36178 76432 36184
rect 76196 36168 76248 36174
rect 76196 36110 76248 36116
rect 76288 36168 76340 36174
rect 76288 36110 76340 36116
rect 75828 36032 75880 36038
rect 75828 35974 75880 35980
rect 75840 35698 75868 35974
rect 75828 35692 75880 35698
rect 75828 35634 75880 35640
rect 76208 34678 76236 36110
rect 70308 34672 70360 34678
rect 70308 34614 70360 34620
rect 71320 34672 71372 34678
rect 71320 34614 71372 34620
rect 74080 34672 74132 34678
rect 74080 34614 74132 34620
rect 76196 34672 76248 34678
rect 76196 34614 76248 34620
rect 70124 34536 70176 34542
rect 70124 34478 70176 34484
rect 70320 34202 70348 34614
rect 77484 34604 77536 34610
rect 77484 34546 77536 34552
rect 71872 34536 71924 34542
rect 71872 34478 71924 34484
rect 70308 34196 70360 34202
rect 70308 34138 70360 34144
rect 68008 34060 68060 34066
rect 68008 34002 68060 34008
rect 68928 34060 68980 34066
rect 68928 34002 68980 34008
rect 71884 33998 71912 34478
rect 77496 34105 77524 34546
rect 77482 34096 77538 34105
rect 77482 34031 77538 34040
rect 66904 33992 66956 33998
rect 66904 33934 66956 33940
rect 71872 33992 71924 33998
rect 71872 33934 71924 33940
rect 66260 33856 66312 33862
rect 66260 33798 66312 33804
rect 5794 33756 6102 33765
rect 5794 33754 5800 33756
rect 5856 33754 5880 33756
rect 5936 33754 5960 33756
rect 6016 33754 6040 33756
rect 6096 33754 6102 33756
rect 5856 33702 5858 33754
rect 6038 33702 6040 33754
rect 5794 33700 5800 33702
rect 5856 33700 5880 33702
rect 5936 33700 5960 33702
rect 6016 33700 6040 33702
rect 6096 33700 6102 33702
rect 5794 33691 6102 33700
rect 36514 33756 36822 33765
rect 36514 33754 36520 33756
rect 36576 33754 36600 33756
rect 36656 33754 36680 33756
rect 36736 33754 36760 33756
rect 36816 33754 36822 33756
rect 36576 33702 36578 33754
rect 36758 33702 36760 33754
rect 36514 33700 36520 33702
rect 36576 33700 36600 33702
rect 36656 33700 36680 33702
rect 36736 33700 36760 33702
rect 36816 33700 36822 33702
rect 36514 33691 36822 33700
rect 66272 33522 66300 33798
rect 66916 33658 66944 33934
rect 67234 33756 67542 33765
rect 67234 33754 67240 33756
rect 67296 33754 67320 33756
rect 67376 33754 67400 33756
rect 67456 33754 67480 33756
rect 67536 33754 67542 33756
rect 67296 33702 67298 33754
rect 67478 33702 67480 33754
rect 67234 33700 67240 33702
rect 67296 33700 67320 33702
rect 67376 33700 67400 33702
rect 67456 33700 67480 33702
rect 67536 33700 67542 33702
rect 67234 33691 67542 33700
rect 66904 33652 66956 33658
rect 66904 33594 66956 33600
rect 66260 33516 66312 33522
rect 66260 33458 66312 33464
rect 5134 33212 5442 33221
rect 5134 33210 5140 33212
rect 5196 33210 5220 33212
rect 5276 33210 5300 33212
rect 5356 33210 5380 33212
rect 5436 33210 5442 33212
rect 5196 33158 5198 33210
rect 5378 33158 5380 33210
rect 5134 33156 5140 33158
rect 5196 33156 5220 33158
rect 5276 33156 5300 33158
rect 5356 33156 5380 33158
rect 5436 33156 5442 33158
rect 5134 33147 5442 33156
rect 35854 33212 36162 33221
rect 35854 33210 35860 33212
rect 35916 33210 35940 33212
rect 35996 33210 36020 33212
rect 36076 33210 36100 33212
rect 36156 33210 36162 33212
rect 35916 33158 35918 33210
rect 36098 33158 36100 33210
rect 35854 33156 35860 33158
rect 35916 33156 35940 33158
rect 35996 33156 36020 33158
rect 36076 33156 36100 33158
rect 36156 33156 36162 33158
rect 35854 33147 36162 33156
rect 66574 33212 66882 33221
rect 66574 33210 66580 33212
rect 66636 33210 66660 33212
rect 66716 33210 66740 33212
rect 66796 33210 66820 33212
rect 66876 33210 66882 33212
rect 66636 33158 66638 33210
rect 66818 33158 66820 33210
rect 66574 33156 66580 33158
rect 66636 33156 66660 33158
rect 66716 33156 66740 33158
rect 66796 33156 66820 33158
rect 66876 33156 66882 33158
rect 66574 33147 66882 33156
rect 5794 32668 6102 32677
rect 5794 32666 5800 32668
rect 5856 32666 5880 32668
rect 5936 32666 5960 32668
rect 6016 32666 6040 32668
rect 6096 32666 6102 32668
rect 5856 32614 5858 32666
rect 6038 32614 6040 32666
rect 5794 32612 5800 32614
rect 5856 32612 5880 32614
rect 5936 32612 5960 32614
rect 6016 32612 6040 32614
rect 6096 32612 6102 32614
rect 5794 32603 6102 32612
rect 36514 32668 36822 32677
rect 36514 32666 36520 32668
rect 36576 32666 36600 32668
rect 36656 32666 36680 32668
rect 36736 32666 36760 32668
rect 36816 32666 36822 32668
rect 36576 32614 36578 32666
rect 36758 32614 36760 32666
rect 36514 32612 36520 32614
rect 36576 32612 36600 32614
rect 36656 32612 36680 32614
rect 36736 32612 36760 32614
rect 36816 32612 36822 32614
rect 36514 32603 36822 32612
rect 67234 32668 67542 32677
rect 67234 32666 67240 32668
rect 67296 32666 67320 32668
rect 67376 32666 67400 32668
rect 67456 32666 67480 32668
rect 67536 32666 67542 32668
rect 67296 32614 67298 32666
rect 67478 32614 67480 32666
rect 67234 32612 67240 32614
rect 67296 32612 67320 32614
rect 67376 32612 67400 32614
rect 67456 32612 67480 32614
rect 67536 32612 67542 32614
rect 67234 32603 67542 32612
rect 1216 32224 1268 32230
rect 1216 32166 1268 32172
rect 1228 32065 1256 32166
rect 5134 32124 5442 32133
rect 5134 32122 5140 32124
rect 5196 32122 5220 32124
rect 5276 32122 5300 32124
rect 5356 32122 5380 32124
rect 5436 32122 5442 32124
rect 5196 32070 5198 32122
rect 5378 32070 5380 32122
rect 5134 32068 5140 32070
rect 5196 32068 5220 32070
rect 5276 32068 5300 32070
rect 5356 32068 5380 32070
rect 5436 32068 5442 32070
rect 1214 32056 1270 32065
rect 5134 32059 5442 32068
rect 35854 32124 36162 32133
rect 35854 32122 35860 32124
rect 35916 32122 35940 32124
rect 35996 32122 36020 32124
rect 36076 32122 36100 32124
rect 36156 32122 36162 32124
rect 35916 32070 35918 32122
rect 36098 32070 36100 32122
rect 35854 32068 35860 32070
rect 35916 32068 35940 32070
rect 35996 32068 36020 32070
rect 36076 32068 36100 32070
rect 36156 32068 36162 32070
rect 35854 32059 36162 32068
rect 66574 32124 66882 32133
rect 66574 32122 66580 32124
rect 66636 32122 66660 32124
rect 66716 32122 66740 32124
rect 66796 32122 66820 32124
rect 66876 32122 66882 32124
rect 66636 32070 66638 32122
rect 66818 32070 66820 32122
rect 66574 32068 66580 32070
rect 66636 32068 66660 32070
rect 66716 32068 66740 32070
rect 66796 32068 66820 32070
rect 66876 32068 66882 32070
rect 66574 32059 66882 32068
rect 1214 31991 1270 32000
rect 5794 31580 6102 31589
rect 5794 31578 5800 31580
rect 5856 31578 5880 31580
rect 5936 31578 5960 31580
rect 6016 31578 6040 31580
rect 6096 31578 6102 31580
rect 5856 31526 5858 31578
rect 6038 31526 6040 31578
rect 5794 31524 5800 31526
rect 5856 31524 5880 31526
rect 5936 31524 5960 31526
rect 6016 31524 6040 31526
rect 6096 31524 6102 31526
rect 5794 31515 6102 31524
rect 36514 31580 36822 31589
rect 36514 31578 36520 31580
rect 36576 31578 36600 31580
rect 36656 31578 36680 31580
rect 36736 31578 36760 31580
rect 36816 31578 36822 31580
rect 36576 31526 36578 31578
rect 36758 31526 36760 31578
rect 36514 31524 36520 31526
rect 36576 31524 36600 31526
rect 36656 31524 36680 31526
rect 36736 31524 36760 31526
rect 36816 31524 36822 31526
rect 36514 31515 36822 31524
rect 67234 31580 67542 31589
rect 67234 31578 67240 31580
rect 67296 31578 67320 31580
rect 67376 31578 67400 31580
rect 67456 31578 67480 31580
rect 67536 31578 67542 31580
rect 67296 31526 67298 31578
rect 67478 31526 67480 31578
rect 67234 31524 67240 31526
rect 67296 31524 67320 31526
rect 67376 31524 67400 31526
rect 67456 31524 67480 31526
rect 67536 31524 67542 31526
rect 67234 31515 67542 31524
rect 5134 31036 5442 31045
rect 5134 31034 5140 31036
rect 5196 31034 5220 31036
rect 5276 31034 5300 31036
rect 5356 31034 5380 31036
rect 5436 31034 5442 31036
rect 5196 30982 5198 31034
rect 5378 30982 5380 31034
rect 5134 30980 5140 30982
rect 5196 30980 5220 30982
rect 5276 30980 5300 30982
rect 5356 30980 5380 30982
rect 5436 30980 5442 30982
rect 5134 30971 5442 30980
rect 35854 31036 36162 31045
rect 35854 31034 35860 31036
rect 35916 31034 35940 31036
rect 35996 31034 36020 31036
rect 36076 31034 36100 31036
rect 36156 31034 36162 31036
rect 35916 30982 35918 31034
rect 36098 30982 36100 31034
rect 35854 30980 35860 30982
rect 35916 30980 35940 30982
rect 35996 30980 36020 30982
rect 36076 30980 36100 30982
rect 36156 30980 36162 30982
rect 35854 30971 36162 30980
rect 66574 31036 66882 31045
rect 66574 31034 66580 31036
rect 66636 31034 66660 31036
rect 66716 31034 66740 31036
rect 66796 31034 66820 31036
rect 66876 31034 66882 31036
rect 66636 30982 66638 31034
rect 66818 30982 66820 31034
rect 66574 30980 66580 30982
rect 66636 30980 66660 30982
rect 66716 30980 66740 30982
rect 66796 30980 66820 30982
rect 66876 30980 66882 30982
rect 66574 30971 66882 30980
rect 5794 30492 6102 30501
rect 5794 30490 5800 30492
rect 5856 30490 5880 30492
rect 5936 30490 5960 30492
rect 6016 30490 6040 30492
rect 6096 30490 6102 30492
rect 5856 30438 5858 30490
rect 6038 30438 6040 30490
rect 5794 30436 5800 30438
rect 5856 30436 5880 30438
rect 5936 30436 5960 30438
rect 6016 30436 6040 30438
rect 6096 30436 6102 30438
rect 5794 30427 6102 30436
rect 36514 30492 36822 30501
rect 36514 30490 36520 30492
rect 36576 30490 36600 30492
rect 36656 30490 36680 30492
rect 36736 30490 36760 30492
rect 36816 30490 36822 30492
rect 36576 30438 36578 30490
rect 36758 30438 36760 30490
rect 36514 30436 36520 30438
rect 36576 30436 36600 30438
rect 36656 30436 36680 30438
rect 36736 30436 36760 30438
rect 36816 30436 36822 30438
rect 36514 30427 36822 30436
rect 67234 30492 67542 30501
rect 67234 30490 67240 30492
rect 67296 30490 67320 30492
rect 67376 30490 67400 30492
rect 67456 30490 67480 30492
rect 67536 30490 67542 30492
rect 67296 30438 67298 30490
rect 67478 30438 67480 30490
rect 67234 30436 67240 30438
rect 67296 30436 67320 30438
rect 67376 30436 67400 30438
rect 67456 30436 67480 30438
rect 67536 30436 67542 30438
rect 67234 30427 67542 30436
rect 5134 29948 5442 29957
rect 5134 29946 5140 29948
rect 5196 29946 5220 29948
rect 5276 29946 5300 29948
rect 5356 29946 5380 29948
rect 5436 29946 5442 29948
rect 5196 29894 5198 29946
rect 5378 29894 5380 29946
rect 5134 29892 5140 29894
rect 5196 29892 5220 29894
rect 5276 29892 5300 29894
rect 5356 29892 5380 29894
rect 5436 29892 5442 29894
rect 5134 29883 5442 29892
rect 35854 29948 36162 29957
rect 35854 29946 35860 29948
rect 35916 29946 35940 29948
rect 35996 29946 36020 29948
rect 36076 29946 36100 29948
rect 36156 29946 36162 29948
rect 35916 29894 35918 29946
rect 36098 29894 36100 29946
rect 35854 29892 35860 29894
rect 35916 29892 35940 29894
rect 35996 29892 36020 29894
rect 36076 29892 36100 29894
rect 36156 29892 36162 29894
rect 35854 29883 36162 29892
rect 66574 29948 66882 29957
rect 66574 29946 66580 29948
rect 66636 29946 66660 29948
rect 66716 29946 66740 29948
rect 66796 29946 66820 29948
rect 66876 29946 66882 29948
rect 66636 29894 66638 29946
rect 66818 29894 66820 29946
rect 66574 29892 66580 29894
rect 66636 29892 66660 29894
rect 66716 29892 66740 29894
rect 66796 29892 66820 29894
rect 66876 29892 66882 29894
rect 66574 29883 66882 29892
rect 5794 29404 6102 29413
rect 5794 29402 5800 29404
rect 5856 29402 5880 29404
rect 5936 29402 5960 29404
rect 6016 29402 6040 29404
rect 6096 29402 6102 29404
rect 5856 29350 5858 29402
rect 6038 29350 6040 29402
rect 5794 29348 5800 29350
rect 5856 29348 5880 29350
rect 5936 29348 5960 29350
rect 6016 29348 6040 29350
rect 6096 29348 6102 29350
rect 5794 29339 6102 29348
rect 36514 29404 36822 29413
rect 36514 29402 36520 29404
rect 36576 29402 36600 29404
rect 36656 29402 36680 29404
rect 36736 29402 36760 29404
rect 36816 29402 36822 29404
rect 36576 29350 36578 29402
rect 36758 29350 36760 29402
rect 36514 29348 36520 29350
rect 36576 29348 36600 29350
rect 36656 29348 36680 29350
rect 36736 29348 36760 29350
rect 36816 29348 36822 29350
rect 36514 29339 36822 29348
rect 67234 29404 67542 29413
rect 67234 29402 67240 29404
rect 67296 29402 67320 29404
rect 67376 29402 67400 29404
rect 67456 29402 67480 29404
rect 67536 29402 67542 29404
rect 67296 29350 67298 29402
rect 67478 29350 67480 29402
rect 67234 29348 67240 29350
rect 67296 29348 67320 29350
rect 67376 29348 67400 29350
rect 67456 29348 67480 29350
rect 67536 29348 67542 29350
rect 67234 29339 67542 29348
rect 2320 29028 2372 29034
rect 2320 28970 2372 28976
rect 2332 28665 2360 28970
rect 5134 28860 5442 28869
rect 5134 28858 5140 28860
rect 5196 28858 5220 28860
rect 5276 28858 5300 28860
rect 5356 28858 5380 28860
rect 5436 28858 5442 28860
rect 5196 28806 5198 28858
rect 5378 28806 5380 28858
rect 5134 28804 5140 28806
rect 5196 28804 5220 28806
rect 5276 28804 5300 28806
rect 5356 28804 5380 28806
rect 5436 28804 5442 28806
rect 5134 28795 5442 28804
rect 35854 28860 36162 28869
rect 35854 28858 35860 28860
rect 35916 28858 35940 28860
rect 35996 28858 36020 28860
rect 36076 28858 36100 28860
rect 36156 28858 36162 28860
rect 35916 28806 35918 28858
rect 36098 28806 36100 28858
rect 35854 28804 35860 28806
rect 35916 28804 35940 28806
rect 35996 28804 36020 28806
rect 36076 28804 36100 28806
rect 36156 28804 36162 28806
rect 35854 28795 36162 28804
rect 66574 28860 66882 28869
rect 66574 28858 66580 28860
rect 66636 28858 66660 28860
rect 66716 28858 66740 28860
rect 66796 28858 66820 28860
rect 66876 28858 66882 28860
rect 66636 28806 66638 28858
rect 66818 28806 66820 28858
rect 66574 28804 66580 28806
rect 66636 28804 66660 28806
rect 66716 28804 66740 28806
rect 66796 28804 66820 28806
rect 66876 28804 66882 28806
rect 66574 28795 66882 28804
rect 2318 28656 2374 28665
rect 2318 28591 2374 28600
rect 5794 28316 6102 28325
rect 5794 28314 5800 28316
rect 5856 28314 5880 28316
rect 5936 28314 5960 28316
rect 6016 28314 6040 28316
rect 6096 28314 6102 28316
rect 5856 28262 5858 28314
rect 6038 28262 6040 28314
rect 5794 28260 5800 28262
rect 5856 28260 5880 28262
rect 5936 28260 5960 28262
rect 6016 28260 6040 28262
rect 6096 28260 6102 28262
rect 5794 28251 6102 28260
rect 36514 28316 36822 28325
rect 36514 28314 36520 28316
rect 36576 28314 36600 28316
rect 36656 28314 36680 28316
rect 36736 28314 36760 28316
rect 36816 28314 36822 28316
rect 36576 28262 36578 28314
rect 36758 28262 36760 28314
rect 36514 28260 36520 28262
rect 36576 28260 36600 28262
rect 36656 28260 36680 28262
rect 36736 28260 36760 28262
rect 36816 28260 36822 28262
rect 36514 28251 36822 28260
rect 67234 28316 67542 28325
rect 67234 28314 67240 28316
rect 67296 28314 67320 28316
rect 67376 28314 67400 28316
rect 67456 28314 67480 28316
rect 67536 28314 67542 28316
rect 67296 28262 67298 28314
rect 67478 28262 67480 28314
rect 67234 28260 67240 28262
rect 67296 28260 67320 28262
rect 67376 28260 67400 28262
rect 67456 28260 67480 28262
rect 67536 28260 67542 28262
rect 67234 28251 67542 28260
rect 1216 28008 1268 28014
rect 1214 27976 1216 27985
rect 1268 27976 1270 27985
rect 1214 27911 1270 27920
rect 5134 27772 5442 27781
rect 5134 27770 5140 27772
rect 5196 27770 5220 27772
rect 5276 27770 5300 27772
rect 5356 27770 5380 27772
rect 5436 27770 5442 27772
rect 5196 27718 5198 27770
rect 5378 27718 5380 27770
rect 5134 27716 5140 27718
rect 5196 27716 5220 27718
rect 5276 27716 5300 27718
rect 5356 27716 5380 27718
rect 5436 27716 5442 27718
rect 5134 27707 5442 27716
rect 35854 27772 36162 27781
rect 35854 27770 35860 27772
rect 35916 27770 35940 27772
rect 35996 27770 36020 27772
rect 36076 27770 36100 27772
rect 36156 27770 36162 27772
rect 35916 27718 35918 27770
rect 36098 27718 36100 27770
rect 35854 27716 35860 27718
rect 35916 27716 35940 27718
rect 35996 27716 36020 27718
rect 36076 27716 36100 27718
rect 36156 27716 36162 27718
rect 35854 27707 36162 27716
rect 66574 27772 66882 27781
rect 66574 27770 66580 27772
rect 66636 27770 66660 27772
rect 66716 27770 66740 27772
rect 66796 27770 66820 27772
rect 66876 27770 66882 27772
rect 66636 27718 66638 27770
rect 66818 27718 66820 27770
rect 66574 27716 66580 27718
rect 66636 27716 66660 27718
rect 66716 27716 66740 27718
rect 66796 27716 66820 27718
rect 66876 27716 66882 27718
rect 66574 27707 66882 27716
rect 5794 27228 6102 27237
rect 5794 27226 5800 27228
rect 5856 27226 5880 27228
rect 5936 27226 5960 27228
rect 6016 27226 6040 27228
rect 6096 27226 6102 27228
rect 5856 27174 5858 27226
rect 6038 27174 6040 27226
rect 5794 27172 5800 27174
rect 5856 27172 5880 27174
rect 5936 27172 5960 27174
rect 6016 27172 6040 27174
rect 6096 27172 6102 27174
rect 5794 27163 6102 27172
rect 36514 27228 36822 27237
rect 36514 27226 36520 27228
rect 36576 27226 36600 27228
rect 36656 27226 36680 27228
rect 36736 27226 36760 27228
rect 36816 27226 36822 27228
rect 36576 27174 36578 27226
rect 36758 27174 36760 27226
rect 36514 27172 36520 27174
rect 36576 27172 36600 27174
rect 36656 27172 36680 27174
rect 36736 27172 36760 27174
rect 36816 27172 36822 27174
rect 36514 27163 36822 27172
rect 67234 27228 67542 27237
rect 67234 27226 67240 27228
rect 67296 27226 67320 27228
rect 67376 27226 67400 27228
rect 67456 27226 67480 27228
rect 67536 27226 67542 27228
rect 67296 27174 67298 27226
rect 67478 27174 67480 27226
rect 67234 27172 67240 27174
rect 67296 27172 67320 27174
rect 67376 27172 67400 27174
rect 67456 27172 67480 27174
rect 67536 27172 67542 27174
rect 67234 27163 67542 27172
rect 1216 26784 1268 26790
rect 1216 26726 1268 26732
rect 1228 26625 1256 26726
rect 5134 26684 5442 26693
rect 5134 26682 5140 26684
rect 5196 26682 5220 26684
rect 5276 26682 5300 26684
rect 5356 26682 5380 26684
rect 5436 26682 5442 26684
rect 5196 26630 5198 26682
rect 5378 26630 5380 26682
rect 5134 26628 5140 26630
rect 5196 26628 5220 26630
rect 5276 26628 5300 26630
rect 5356 26628 5380 26630
rect 5436 26628 5442 26630
rect 1214 26616 1270 26625
rect 5134 26619 5442 26628
rect 35854 26684 36162 26693
rect 35854 26682 35860 26684
rect 35916 26682 35940 26684
rect 35996 26682 36020 26684
rect 36076 26682 36100 26684
rect 36156 26682 36162 26684
rect 35916 26630 35918 26682
rect 36098 26630 36100 26682
rect 35854 26628 35860 26630
rect 35916 26628 35940 26630
rect 35996 26628 36020 26630
rect 36076 26628 36100 26630
rect 36156 26628 36162 26630
rect 35854 26619 36162 26628
rect 66574 26684 66882 26693
rect 66574 26682 66580 26684
rect 66636 26682 66660 26684
rect 66716 26682 66740 26684
rect 66796 26682 66820 26684
rect 66876 26682 66882 26684
rect 66636 26630 66638 26682
rect 66818 26630 66820 26682
rect 66574 26628 66580 26630
rect 66636 26628 66660 26630
rect 66716 26628 66740 26630
rect 66796 26628 66820 26630
rect 66876 26628 66882 26630
rect 66574 26619 66882 26628
rect 1214 26551 1270 26560
rect 2320 26376 2372 26382
rect 2320 26318 2372 26324
rect 2332 25945 2360 26318
rect 5794 26140 6102 26149
rect 5794 26138 5800 26140
rect 5856 26138 5880 26140
rect 5936 26138 5960 26140
rect 6016 26138 6040 26140
rect 6096 26138 6102 26140
rect 5856 26086 5858 26138
rect 6038 26086 6040 26138
rect 5794 26084 5800 26086
rect 5856 26084 5880 26086
rect 5936 26084 5960 26086
rect 6016 26084 6040 26086
rect 6096 26084 6102 26086
rect 5794 26075 6102 26084
rect 36514 26140 36822 26149
rect 36514 26138 36520 26140
rect 36576 26138 36600 26140
rect 36656 26138 36680 26140
rect 36736 26138 36760 26140
rect 36816 26138 36822 26140
rect 36576 26086 36578 26138
rect 36758 26086 36760 26138
rect 36514 26084 36520 26086
rect 36576 26084 36600 26086
rect 36656 26084 36680 26086
rect 36736 26084 36760 26086
rect 36816 26084 36822 26086
rect 36514 26075 36822 26084
rect 67234 26140 67542 26149
rect 67234 26138 67240 26140
rect 67296 26138 67320 26140
rect 67376 26138 67400 26140
rect 67456 26138 67480 26140
rect 67536 26138 67542 26140
rect 67296 26086 67298 26138
rect 67478 26086 67480 26138
rect 67234 26084 67240 26086
rect 67296 26084 67320 26086
rect 67376 26084 67400 26086
rect 67456 26084 67480 26086
rect 67536 26084 67542 26086
rect 67234 26075 67542 26084
rect 2318 25936 2374 25945
rect 2318 25871 2374 25880
rect 5134 25596 5442 25605
rect 5134 25594 5140 25596
rect 5196 25594 5220 25596
rect 5276 25594 5300 25596
rect 5356 25594 5380 25596
rect 5436 25594 5442 25596
rect 5196 25542 5198 25594
rect 5378 25542 5380 25594
rect 5134 25540 5140 25542
rect 5196 25540 5220 25542
rect 5276 25540 5300 25542
rect 5356 25540 5380 25542
rect 5436 25540 5442 25542
rect 5134 25531 5442 25540
rect 35854 25596 36162 25605
rect 35854 25594 35860 25596
rect 35916 25594 35940 25596
rect 35996 25594 36020 25596
rect 36076 25594 36100 25596
rect 36156 25594 36162 25596
rect 35916 25542 35918 25594
rect 36098 25542 36100 25594
rect 35854 25540 35860 25542
rect 35916 25540 35940 25542
rect 35996 25540 36020 25542
rect 36076 25540 36100 25542
rect 36156 25540 36162 25542
rect 35854 25531 36162 25540
rect 66574 25596 66882 25605
rect 66574 25594 66580 25596
rect 66636 25594 66660 25596
rect 66716 25594 66740 25596
rect 66796 25594 66820 25596
rect 66876 25594 66882 25596
rect 66636 25542 66638 25594
rect 66818 25542 66820 25594
rect 66574 25540 66580 25542
rect 66636 25540 66660 25542
rect 66716 25540 66740 25542
rect 66796 25540 66820 25542
rect 66876 25540 66882 25542
rect 66574 25531 66882 25540
rect 5794 25052 6102 25061
rect 5794 25050 5800 25052
rect 5856 25050 5880 25052
rect 5936 25050 5960 25052
rect 6016 25050 6040 25052
rect 6096 25050 6102 25052
rect 5856 24998 5858 25050
rect 6038 24998 6040 25050
rect 5794 24996 5800 24998
rect 5856 24996 5880 24998
rect 5936 24996 5960 24998
rect 6016 24996 6040 24998
rect 6096 24996 6102 24998
rect 5794 24987 6102 24996
rect 36514 25052 36822 25061
rect 36514 25050 36520 25052
rect 36576 25050 36600 25052
rect 36656 25050 36680 25052
rect 36736 25050 36760 25052
rect 36816 25050 36822 25052
rect 36576 24998 36578 25050
rect 36758 24998 36760 25050
rect 36514 24996 36520 24998
rect 36576 24996 36600 24998
rect 36656 24996 36680 24998
rect 36736 24996 36760 24998
rect 36816 24996 36822 24998
rect 36514 24987 36822 24996
rect 67234 25052 67542 25061
rect 67234 25050 67240 25052
rect 67296 25050 67320 25052
rect 67376 25050 67400 25052
rect 67456 25050 67480 25052
rect 67536 25050 67542 25052
rect 67296 24998 67298 25050
rect 67478 24998 67480 25050
rect 67234 24996 67240 24998
rect 67296 24996 67320 24998
rect 67376 24996 67400 24998
rect 67456 24996 67480 24998
rect 67536 24996 67542 24998
rect 67234 24987 67542 24996
rect 5134 24508 5442 24517
rect 5134 24506 5140 24508
rect 5196 24506 5220 24508
rect 5276 24506 5300 24508
rect 5356 24506 5380 24508
rect 5436 24506 5442 24508
rect 5196 24454 5198 24506
rect 5378 24454 5380 24506
rect 5134 24452 5140 24454
rect 5196 24452 5220 24454
rect 5276 24452 5300 24454
rect 5356 24452 5380 24454
rect 5436 24452 5442 24454
rect 5134 24443 5442 24452
rect 35854 24508 36162 24517
rect 35854 24506 35860 24508
rect 35916 24506 35940 24508
rect 35996 24506 36020 24508
rect 36076 24506 36100 24508
rect 36156 24506 36162 24508
rect 35916 24454 35918 24506
rect 36098 24454 36100 24506
rect 35854 24452 35860 24454
rect 35916 24452 35940 24454
rect 35996 24452 36020 24454
rect 36076 24452 36100 24454
rect 36156 24452 36162 24454
rect 35854 24443 36162 24452
rect 66574 24508 66882 24517
rect 66574 24506 66580 24508
rect 66636 24506 66660 24508
rect 66716 24506 66740 24508
rect 66796 24506 66820 24508
rect 66876 24506 66882 24508
rect 66636 24454 66638 24506
rect 66818 24454 66820 24506
rect 66574 24452 66580 24454
rect 66636 24452 66660 24454
rect 66716 24452 66740 24454
rect 66796 24452 66820 24454
rect 66876 24452 66882 24454
rect 66574 24443 66882 24452
rect 5794 23964 6102 23973
rect 5794 23962 5800 23964
rect 5856 23962 5880 23964
rect 5936 23962 5960 23964
rect 6016 23962 6040 23964
rect 6096 23962 6102 23964
rect 5856 23910 5858 23962
rect 6038 23910 6040 23962
rect 5794 23908 5800 23910
rect 5856 23908 5880 23910
rect 5936 23908 5960 23910
rect 6016 23908 6040 23910
rect 6096 23908 6102 23910
rect 5794 23899 6102 23908
rect 36514 23964 36822 23973
rect 36514 23962 36520 23964
rect 36576 23962 36600 23964
rect 36656 23962 36680 23964
rect 36736 23962 36760 23964
rect 36816 23962 36822 23964
rect 36576 23910 36578 23962
rect 36758 23910 36760 23962
rect 36514 23908 36520 23910
rect 36576 23908 36600 23910
rect 36656 23908 36680 23910
rect 36736 23908 36760 23910
rect 36816 23908 36822 23910
rect 36514 23899 36822 23908
rect 67234 23964 67542 23973
rect 67234 23962 67240 23964
rect 67296 23962 67320 23964
rect 67376 23962 67400 23964
rect 67456 23962 67480 23964
rect 67536 23962 67542 23964
rect 67296 23910 67298 23962
rect 67478 23910 67480 23962
rect 67234 23908 67240 23910
rect 67296 23908 67320 23910
rect 67376 23908 67400 23910
rect 67456 23908 67480 23910
rect 67536 23908 67542 23910
rect 67234 23899 67542 23908
rect 2320 23520 2372 23526
rect 2320 23462 2372 23468
rect 2332 23225 2360 23462
rect 5134 23420 5442 23429
rect 5134 23418 5140 23420
rect 5196 23418 5220 23420
rect 5276 23418 5300 23420
rect 5356 23418 5380 23420
rect 5436 23418 5442 23420
rect 5196 23366 5198 23418
rect 5378 23366 5380 23418
rect 5134 23364 5140 23366
rect 5196 23364 5220 23366
rect 5276 23364 5300 23366
rect 5356 23364 5380 23366
rect 5436 23364 5442 23366
rect 5134 23355 5442 23364
rect 35854 23420 36162 23429
rect 35854 23418 35860 23420
rect 35916 23418 35940 23420
rect 35996 23418 36020 23420
rect 36076 23418 36100 23420
rect 36156 23418 36162 23420
rect 35916 23366 35918 23418
rect 36098 23366 36100 23418
rect 35854 23364 35860 23366
rect 35916 23364 35940 23366
rect 35996 23364 36020 23366
rect 36076 23364 36100 23366
rect 36156 23364 36162 23366
rect 35854 23355 36162 23364
rect 66574 23420 66882 23429
rect 66574 23418 66580 23420
rect 66636 23418 66660 23420
rect 66716 23418 66740 23420
rect 66796 23418 66820 23420
rect 66876 23418 66882 23420
rect 66636 23366 66638 23418
rect 66818 23366 66820 23418
rect 66574 23364 66580 23366
rect 66636 23364 66660 23366
rect 66716 23364 66740 23366
rect 66796 23364 66820 23366
rect 66876 23364 66882 23366
rect 66574 23355 66882 23364
rect 2318 23216 2374 23225
rect 2318 23151 2374 23160
rect 5794 22876 6102 22885
rect 5794 22874 5800 22876
rect 5856 22874 5880 22876
rect 5936 22874 5960 22876
rect 6016 22874 6040 22876
rect 6096 22874 6102 22876
rect 5856 22822 5858 22874
rect 6038 22822 6040 22874
rect 5794 22820 5800 22822
rect 5856 22820 5880 22822
rect 5936 22820 5960 22822
rect 6016 22820 6040 22822
rect 6096 22820 6102 22822
rect 5794 22811 6102 22820
rect 36514 22876 36822 22885
rect 36514 22874 36520 22876
rect 36576 22874 36600 22876
rect 36656 22874 36680 22876
rect 36736 22874 36760 22876
rect 36816 22874 36822 22876
rect 36576 22822 36578 22874
rect 36758 22822 36760 22874
rect 36514 22820 36520 22822
rect 36576 22820 36600 22822
rect 36656 22820 36680 22822
rect 36736 22820 36760 22822
rect 36816 22820 36822 22822
rect 36514 22811 36822 22820
rect 67234 22876 67542 22885
rect 67234 22874 67240 22876
rect 67296 22874 67320 22876
rect 67376 22874 67400 22876
rect 67456 22874 67480 22876
rect 67536 22874 67542 22876
rect 67296 22822 67298 22874
rect 67478 22822 67480 22874
rect 67234 22820 67240 22822
rect 67296 22820 67320 22822
rect 67376 22820 67400 22822
rect 67456 22820 67480 22822
rect 67536 22820 67542 22822
rect 67234 22811 67542 22820
rect 5134 22332 5442 22341
rect 5134 22330 5140 22332
rect 5196 22330 5220 22332
rect 5276 22330 5300 22332
rect 5356 22330 5380 22332
rect 5436 22330 5442 22332
rect 5196 22278 5198 22330
rect 5378 22278 5380 22330
rect 5134 22276 5140 22278
rect 5196 22276 5220 22278
rect 5276 22276 5300 22278
rect 5356 22276 5380 22278
rect 5436 22276 5442 22278
rect 5134 22267 5442 22276
rect 35854 22332 36162 22341
rect 35854 22330 35860 22332
rect 35916 22330 35940 22332
rect 35996 22330 36020 22332
rect 36076 22330 36100 22332
rect 36156 22330 36162 22332
rect 35916 22278 35918 22330
rect 36098 22278 36100 22330
rect 35854 22276 35860 22278
rect 35916 22276 35940 22278
rect 35996 22276 36020 22278
rect 36076 22276 36100 22278
rect 36156 22276 36162 22278
rect 35854 22267 36162 22276
rect 66574 22332 66882 22341
rect 66574 22330 66580 22332
rect 66636 22330 66660 22332
rect 66716 22330 66740 22332
rect 66796 22330 66820 22332
rect 66876 22330 66882 22332
rect 66636 22278 66638 22330
rect 66818 22278 66820 22330
rect 66574 22276 66580 22278
rect 66636 22276 66660 22278
rect 66716 22276 66740 22278
rect 66796 22276 66820 22278
rect 66876 22276 66882 22278
rect 66574 22267 66882 22276
rect 5794 21788 6102 21797
rect 5794 21786 5800 21788
rect 5856 21786 5880 21788
rect 5936 21786 5960 21788
rect 6016 21786 6040 21788
rect 6096 21786 6102 21788
rect 5856 21734 5858 21786
rect 6038 21734 6040 21786
rect 5794 21732 5800 21734
rect 5856 21732 5880 21734
rect 5936 21732 5960 21734
rect 6016 21732 6040 21734
rect 6096 21732 6102 21734
rect 5794 21723 6102 21732
rect 36514 21788 36822 21797
rect 36514 21786 36520 21788
rect 36576 21786 36600 21788
rect 36656 21786 36680 21788
rect 36736 21786 36760 21788
rect 36816 21786 36822 21788
rect 36576 21734 36578 21786
rect 36758 21734 36760 21786
rect 36514 21732 36520 21734
rect 36576 21732 36600 21734
rect 36656 21732 36680 21734
rect 36736 21732 36760 21734
rect 36816 21732 36822 21734
rect 36514 21723 36822 21732
rect 67234 21788 67542 21797
rect 67234 21786 67240 21788
rect 67296 21786 67320 21788
rect 67376 21786 67400 21788
rect 67456 21786 67480 21788
rect 67536 21786 67542 21788
rect 67296 21734 67298 21786
rect 67478 21734 67480 21786
rect 67234 21732 67240 21734
rect 67296 21732 67320 21734
rect 67376 21732 67400 21734
rect 67456 21732 67480 21734
rect 67536 21732 67542 21734
rect 67234 21723 67542 21732
rect 77576 21344 77628 21350
rect 77576 21286 77628 21292
rect 5134 21244 5442 21253
rect 5134 21242 5140 21244
rect 5196 21242 5220 21244
rect 5276 21242 5300 21244
rect 5356 21242 5380 21244
rect 5436 21242 5442 21244
rect 5196 21190 5198 21242
rect 5378 21190 5380 21242
rect 5134 21188 5140 21190
rect 5196 21188 5220 21190
rect 5276 21188 5300 21190
rect 5356 21188 5380 21190
rect 5436 21188 5442 21190
rect 5134 21179 5442 21188
rect 35854 21244 36162 21253
rect 35854 21242 35860 21244
rect 35916 21242 35940 21244
rect 35996 21242 36020 21244
rect 36076 21242 36100 21244
rect 36156 21242 36162 21244
rect 35916 21190 35918 21242
rect 36098 21190 36100 21242
rect 35854 21188 35860 21190
rect 35916 21188 35940 21190
rect 35996 21188 36020 21190
rect 36076 21188 36100 21190
rect 36156 21188 36162 21190
rect 35854 21179 36162 21188
rect 66574 21244 66882 21253
rect 66574 21242 66580 21244
rect 66636 21242 66660 21244
rect 66716 21242 66740 21244
rect 66796 21242 66820 21244
rect 66876 21242 66882 21244
rect 66636 21190 66638 21242
rect 66818 21190 66820 21242
rect 66574 21188 66580 21190
rect 66636 21188 66660 21190
rect 66716 21188 66740 21190
rect 66796 21188 66820 21190
rect 66876 21188 66882 21190
rect 66574 21179 66882 21188
rect 77588 21185 77616 21286
rect 77574 21176 77630 21185
rect 77574 21111 77630 21120
rect 5794 20700 6102 20709
rect 5794 20698 5800 20700
rect 5856 20698 5880 20700
rect 5936 20698 5960 20700
rect 6016 20698 6040 20700
rect 6096 20698 6102 20700
rect 5856 20646 5858 20698
rect 6038 20646 6040 20698
rect 5794 20644 5800 20646
rect 5856 20644 5880 20646
rect 5936 20644 5960 20646
rect 6016 20644 6040 20646
rect 6096 20644 6102 20646
rect 5794 20635 6102 20644
rect 36514 20700 36822 20709
rect 36514 20698 36520 20700
rect 36576 20698 36600 20700
rect 36656 20698 36680 20700
rect 36736 20698 36760 20700
rect 36816 20698 36822 20700
rect 36576 20646 36578 20698
rect 36758 20646 36760 20698
rect 36514 20644 36520 20646
rect 36576 20644 36600 20646
rect 36656 20644 36680 20646
rect 36736 20644 36760 20646
rect 36816 20644 36822 20646
rect 36514 20635 36822 20644
rect 67234 20700 67542 20709
rect 67234 20698 67240 20700
rect 67296 20698 67320 20700
rect 67376 20698 67400 20700
rect 67456 20698 67480 20700
rect 67536 20698 67542 20700
rect 67296 20646 67298 20698
rect 67478 20646 67480 20698
rect 67234 20644 67240 20646
rect 67296 20644 67320 20646
rect 67376 20644 67400 20646
rect 67456 20644 67480 20646
rect 67536 20644 67542 20646
rect 67234 20635 67542 20644
rect 5134 20156 5442 20165
rect 5134 20154 5140 20156
rect 5196 20154 5220 20156
rect 5276 20154 5300 20156
rect 5356 20154 5380 20156
rect 5436 20154 5442 20156
rect 5196 20102 5198 20154
rect 5378 20102 5380 20154
rect 5134 20100 5140 20102
rect 5196 20100 5220 20102
rect 5276 20100 5300 20102
rect 5356 20100 5380 20102
rect 5436 20100 5442 20102
rect 5134 20091 5442 20100
rect 35854 20156 36162 20165
rect 35854 20154 35860 20156
rect 35916 20154 35940 20156
rect 35996 20154 36020 20156
rect 36076 20154 36100 20156
rect 36156 20154 36162 20156
rect 35916 20102 35918 20154
rect 36098 20102 36100 20154
rect 35854 20100 35860 20102
rect 35916 20100 35940 20102
rect 35996 20100 36020 20102
rect 36076 20100 36100 20102
rect 36156 20100 36162 20102
rect 35854 20091 36162 20100
rect 66574 20156 66882 20165
rect 66574 20154 66580 20156
rect 66636 20154 66660 20156
rect 66716 20154 66740 20156
rect 66796 20154 66820 20156
rect 66876 20154 66882 20156
rect 66636 20102 66638 20154
rect 66818 20102 66820 20154
rect 66574 20100 66580 20102
rect 66636 20100 66660 20102
rect 66716 20100 66740 20102
rect 66796 20100 66820 20102
rect 66876 20100 66882 20102
rect 66574 20091 66882 20100
rect 5794 19612 6102 19621
rect 5794 19610 5800 19612
rect 5856 19610 5880 19612
rect 5936 19610 5960 19612
rect 6016 19610 6040 19612
rect 6096 19610 6102 19612
rect 5856 19558 5858 19610
rect 6038 19558 6040 19610
rect 5794 19556 5800 19558
rect 5856 19556 5880 19558
rect 5936 19556 5960 19558
rect 6016 19556 6040 19558
rect 6096 19556 6102 19558
rect 5794 19547 6102 19556
rect 36514 19612 36822 19621
rect 36514 19610 36520 19612
rect 36576 19610 36600 19612
rect 36656 19610 36680 19612
rect 36736 19610 36760 19612
rect 36816 19610 36822 19612
rect 36576 19558 36578 19610
rect 36758 19558 36760 19610
rect 36514 19556 36520 19558
rect 36576 19556 36600 19558
rect 36656 19556 36680 19558
rect 36736 19556 36760 19558
rect 36816 19556 36822 19558
rect 36514 19547 36822 19556
rect 67234 19612 67542 19621
rect 67234 19610 67240 19612
rect 67296 19610 67320 19612
rect 67376 19610 67400 19612
rect 67456 19610 67480 19612
rect 67536 19610 67542 19612
rect 67296 19558 67298 19610
rect 67478 19558 67480 19610
rect 67234 19556 67240 19558
rect 67296 19556 67320 19558
rect 67376 19556 67400 19558
rect 67456 19556 67480 19558
rect 67536 19556 67542 19558
rect 67234 19547 67542 19556
rect 5134 19068 5442 19077
rect 5134 19066 5140 19068
rect 5196 19066 5220 19068
rect 5276 19066 5300 19068
rect 5356 19066 5380 19068
rect 5436 19066 5442 19068
rect 5196 19014 5198 19066
rect 5378 19014 5380 19066
rect 5134 19012 5140 19014
rect 5196 19012 5220 19014
rect 5276 19012 5300 19014
rect 5356 19012 5380 19014
rect 5436 19012 5442 19014
rect 5134 19003 5442 19012
rect 35854 19068 36162 19077
rect 35854 19066 35860 19068
rect 35916 19066 35940 19068
rect 35996 19066 36020 19068
rect 36076 19066 36100 19068
rect 36156 19066 36162 19068
rect 35916 19014 35918 19066
rect 36098 19014 36100 19066
rect 35854 19012 35860 19014
rect 35916 19012 35940 19014
rect 35996 19012 36020 19014
rect 36076 19012 36100 19014
rect 36156 19012 36162 19014
rect 35854 19003 36162 19012
rect 66574 19068 66882 19077
rect 66574 19066 66580 19068
rect 66636 19066 66660 19068
rect 66716 19066 66740 19068
rect 66796 19066 66820 19068
rect 66876 19066 66882 19068
rect 66636 19014 66638 19066
rect 66818 19014 66820 19066
rect 66574 19012 66580 19014
rect 66636 19012 66660 19014
rect 66716 19012 66740 19014
rect 66796 19012 66820 19014
rect 66876 19012 66882 19014
rect 66574 19003 66882 19012
rect 5794 18524 6102 18533
rect 5794 18522 5800 18524
rect 5856 18522 5880 18524
rect 5936 18522 5960 18524
rect 6016 18522 6040 18524
rect 6096 18522 6102 18524
rect 5856 18470 5858 18522
rect 6038 18470 6040 18522
rect 5794 18468 5800 18470
rect 5856 18468 5880 18470
rect 5936 18468 5960 18470
rect 6016 18468 6040 18470
rect 6096 18468 6102 18470
rect 5794 18459 6102 18468
rect 36514 18524 36822 18533
rect 36514 18522 36520 18524
rect 36576 18522 36600 18524
rect 36656 18522 36680 18524
rect 36736 18522 36760 18524
rect 36816 18522 36822 18524
rect 36576 18470 36578 18522
rect 36758 18470 36760 18522
rect 36514 18468 36520 18470
rect 36576 18468 36600 18470
rect 36656 18468 36680 18470
rect 36736 18468 36760 18470
rect 36816 18468 36822 18470
rect 36514 18459 36822 18468
rect 67234 18524 67542 18533
rect 67234 18522 67240 18524
rect 67296 18522 67320 18524
rect 67376 18522 67400 18524
rect 67456 18522 67480 18524
rect 67536 18522 67542 18524
rect 67296 18470 67298 18522
rect 67478 18470 67480 18522
rect 67234 18468 67240 18470
rect 67296 18468 67320 18470
rect 67376 18468 67400 18470
rect 67456 18468 67480 18470
rect 67536 18468 67542 18470
rect 67234 18459 67542 18468
rect 5134 17980 5442 17989
rect 5134 17978 5140 17980
rect 5196 17978 5220 17980
rect 5276 17978 5300 17980
rect 5356 17978 5380 17980
rect 5436 17978 5442 17980
rect 5196 17926 5198 17978
rect 5378 17926 5380 17978
rect 5134 17924 5140 17926
rect 5196 17924 5220 17926
rect 5276 17924 5300 17926
rect 5356 17924 5380 17926
rect 5436 17924 5442 17926
rect 5134 17915 5442 17924
rect 35854 17980 36162 17989
rect 35854 17978 35860 17980
rect 35916 17978 35940 17980
rect 35996 17978 36020 17980
rect 36076 17978 36100 17980
rect 36156 17978 36162 17980
rect 35916 17926 35918 17978
rect 36098 17926 36100 17978
rect 35854 17924 35860 17926
rect 35916 17924 35940 17926
rect 35996 17924 36020 17926
rect 36076 17924 36100 17926
rect 36156 17924 36162 17926
rect 35854 17915 36162 17924
rect 66574 17980 66882 17989
rect 66574 17978 66580 17980
rect 66636 17978 66660 17980
rect 66716 17978 66740 17980
rect 66796 17978 66820 17980
rect 66876 17978 66882 17980
rect 66636 17926 66638 17978
rect 66818 17926 66820 17978
rect 66574 17924 66580 17926
rect 66636 17924 66660 17926
rect 66716 17924 66740 17926
rect 66796 17924 66820 17926
rect 66876 17924 66882 17926
rect 66574 17915 66882 17924
rect 5794 17436 6102 17445
rect 5794 17434 5800 17436
rect 5856 17434 5880 17436
rect 5936 17434 5960 17436
rect 6016 17434 6040 17436
rect 6096 17434 6102 17436
rect 5856 17382 5858 17434
rect 6038 17382 6040 17434
rect 5794 17380 5800 17382
rect 5856 17380 5880 17382
rect 5936 17380 5960 17382
rect 6016 17380 6040 17382
rect 6096 17380 6102 17382
rect 5794 17371 6102 17380
rect 36514 17436 36822 17445
rect 36514 17434 36520 17436
rect 36576 17434 36600 17436
rect 36656 17434 36680 17436
rect 36736 17434 36760 17436
rect 36816 17434 36822 17436
rect 36576 17382 36578 17434
rect 36758 17382 36760 17434
rect 36514 17380 36520 17382
rect 36576 17380 36600 17382
rect 36656 17380 36680 17382
rect 36736 17380 36760 17382
rect 36816 17380 36822 17382
rect 36514 17371 36822 17380
rect 67234 17436 67542 17445
rect 67234 17434 67240 17436
rect 67296 17434 67320 17436
rect 67376 17434 67400 17436
rect 67456 17434 67480 17436
rect 67536 17434 67542 17436
rect 67296 17382 67298 17434
rect 67478 17382 67480 17434
rect 67234 17380 67240 17382
rect 67296 17380 67320 17382
rect 67376 17380 67400 17382
rect 67456 17380 67480 17382
rect 67536 17380 67542 17382
rect 67234 17371 67542 17380
rect 5134 16892 5442 16901
rect 5134 16890 5140 16892
rect 5196 16890 5220 16892
rect 5276 16890 5300 16892
rect 5356 16890 5380 16892
rect 5436 16890 5442 16892
rect 5196 16838 5198 16890
rect 5378 16838 5380 16890
rect 5134 16836 5140 16838
rect 5196 16836 5220 16838
rect 5276 16836 5300 16838
rect 5356 16836 5380 16838
rect 5436 16836 5442 16838
rect 5134 16827 5442 16836
rect 35854 16892 36162 16901
rect 35854 16890 35860 16892
rect 35916 16890 35940 16892
rect 35996 16890 36020 16892
rect 36076 16890 36100 16892
rect 36156 16890 36162 16892
rect 35916 16838 35918 16890
rect 36098 16838 36100 16890
rect 35854 16836 35860 16838
rect 35916 16836 35940 16838
rect 35996 16836 36020 16838
rect 36076 16836 36100 16838
rect 36156 16836 36162 16838
rect 35854 16827 36162 16836
rect 66574 16892 66882 16901
rect 66574 16890 66580 16892
rect 66636 16890 66660 16892
rect 66716 16890 66740 16892
rect 66796 16890 66820 16892
rect 66876 16890 66882 16892
rect 66636 16838 66638 16890
rect 66818 16838 66820 16890
rect 66574 16836 66580 16838
rect 66636 16836 66660 16838
rect 66716 16836 66740 16838
rect 66796 16836 66820 16838
rect 66876 16836 66882 16838
rect 66574 16827 66882 16836
rect 77576 16652 77628 16658
rect 77576 16594 77628 16600
rect 77588 16425 77616 16594
rect 77574 16416 77630 16425
rect 5794 16348 6102 16357
rect 5794 16346 5800 16348
rect 5856 16346 5880 16348
rect 5936 16346 5960 16348
rect 6016 16346 6040 16348
rect 6096 16346 6102 16348
rect 5856 16294 5858 16346
rect 6038 16294 6040 16346
rect 5794 16292 5800 16294
rect 5856 16292 5880 16294
rect 5936 16292 5960 16294
rect 6016 16292 6040 16294
rect 6096 16292 6102 16294
rect 5794 16283 6102 16292
rect 36514 16348 36822 16357
rect 36514 16346 36520 16348
rect 36576 16346 36600 16348
rect 36656 16346 36680 16348
rect 36736 16346 36760 16348
rect 36816 16346 36822 16348
rect 36576 16294 36578 16346
rect 36758 16294 36760 16346
rect 36514 16292 36520 16294
rect 36576 16292 36600 16294
rect 36656 16292 36680 16294
rect 36736 16292 36760 16294
rect 36816 16292 36822 16294
rect 36514 16283 36822 16292
rect 67234 16348 67542 16357
rect 77574 16351 77630 16360
rect 67234 16346 67240 16348
rect 67296 16346 67320 16348
rect 67376 16346 67400 16348
rect 67456 16346 67480 16348
rect 67536 16346 67542 16348
rect 67296 16294 67298 16346
rect 67478 16294 67480 16346
rect 67234 16292 67240 16294
rect 67296 16292 67320 16294
rect 67376 16292 67400 16294
rect 67456 16292 67480 16294
rect 67536 16292 67542 16294
rect 67234 16283 67542 16292
rect 5134 15804 5442 15813
rect 5134 15802 5140 15804
rect 5196 15802 5220 15804
rect 5276 15802 5300 15804
rect 5356 15802 5380 15804
rect 5436 15802 5442 15804
rect 5196 15750 5198 15802
rect 5378 15750 5380 15802
rect 5134 15748 5140 15750
rect 5196 15748 5220 15750
rect 5276 15748 5300 15750
rect 5356 15748 5380 15750
rect 5436 15748 5442 15750
rect 5134 15739 5442 15748
rect 35854 15804 36162 15813
rect 35854 15802 35860 15804
rect 35916 15802 35940 15804
rect 35996 15802 36020 15804
rect 36076 15802 36100 15804
rect 36156 15802 36162 15804
rect 35916 15750 35918 15802
rect 36098 15750 36100 15802
rect 35854 15748 35860 15750
rect 35916 15748 35940 15750
rect 35996 15748 36020 15750
rect 36076 15748 36100 15750
rect 36156 15748 36162 15750
rect 35854 15739 36162 15748
rect 66574 15804 66882 15813
rect 66574 15802 66580 15804
rect 66636 15802 66660 15804
rect 66716 15802 66740 15804
rect 66796 15802 66820 15804
rect 66876 15802 66882 15804
rect 66636 15750 66638 15802
rect 66818 15750 66820 15802
rect 66574 15748 66580 15750
rect 66636 15748 66660 15750
rect 66716 15748 66740 15750
rect 66796 15748 66820 15750
rect 66876 15748 66882 15750
rect 66574 15739 66882 15748
rect 5794 15260 6102 15269
rect 5794 15258 5800 15260
rect 5856 15258 5880 15260
rect 5936 15258 5960 15260
rect 6016 15258 6040 15260
rect 6096 15258 6102 15260
rect 5856 15206 5858 15258
rect 6038 15206 6040 15258
rect 5794 15204 5800 15206
rect 5856 15204 5880 15206
rect 5936 15204 5960 15206
rect 6016 15204 6040 15206
rect 6096 15204 6102 15206
rect 5794 15195 6102 15204
rect 36514 15260 36822 15269
rect 36514 15258 36520 15260
rect 36576 15258 36600 15260
rect 36656 15258 36680 15260
rect 36736 15258 36760 15260
rect 36816 15258 36822 15260
rect 36576 15206 36578 15258
rect 36758 15206 36760 15258
rect 36514 15204 36520 15206
rect 36576 15204 36600 15206
rect 36656 15204 36680 15206
rect 36736 15204 36760 15206
rect 36816 15204 36822 15206
rect 36514 15195 36822 15204
rect 67234 15260 67542 15269
rect 67234 15258 67240 15260
rect 67296 15258 67320 15260
rect 67376 15258 67400 15260
rect 67456 15258 67480 15260
rect 67536 15258 67542 15260
rect 67296 15206 67298 15258
rect 67478 15206 67480 15258
rect 67234 15204 67240 15206
rect 67296 15204 67320 15206
rect 67376 15204 67400 15206
rect 67456 15204 67480 15206
rect 67536 15204 67542 15206
rect 67234 15195 67542 15204
rect 5134 14716 5442 14725
rect 5134 14714 5140 14716
rect 5196 14714 5220 14716
rect 5276 14714 5300 14716
rect 5356 14714 5380 14716
rect 5436 14714 5442 14716
rect 5196 14662 5198 14714
rect 5378 14662 5380 14714
rect 5134 14660 5140 14662
rect 5196 14660 5220 14662
rect 5276 14660 5300 14662
rect 5356 14660 5380 14662
rect 5436 14660 5442 14662
rect 5134 14651 5442 14660
rect 35854 14716 36162 14725
rect 35854 14714 35860 14716
rect 35916 14714 35940 14716
rect 35996 14714 36020 14716
rect 36076 14714 36100 14716
rect 36156 14714 36162 14716
rect 35916 14662 35918 14714
rect 36098 14662 36100 14714
rect 35854 14660 35860 14662
rect 35916 14660 35940 14662
rect 35996 14660 36020 14662
rect 36076 14660 36100 14662
rect 36156 14660 36162 14662
rect 35854 14651 36162 14660
rect 66574 14716 66882 14725
rect 66574 14714 66580 14716
rect 66636 14714 66660 14716
rect 66716 14714 66740 14716
rect 66796 14714 66820 14716
rect 66876 14714 66882 14716
rect 66636 14662 66638 14714
rect 66818 14662 66820 14714
rect 66574 14660 66580 14662
rect 66636 14660 66660 14662
rect 66716 14660 66740 14662
rect 66796 14660 66820 14662
rect 66876 14660 66882 14662
rect 66574 14651 66882 14660
rect 5794 14172 6102 14181
rect 5794 14170 5800 14172
rect 5856 14170 5880 14172
rect 5936 14170 5960 14172
rect 6016 14170 6040 14172
rect 6096 14170 6102 14172
rect 5856 14118 5858 14170
rect 6038 14118 6040 14170
rect 5794 14116 5800 14118
rect 5856 14116 5880 14118
rect 5936 14116 5960 14118
rect 6016 14116 6040 14118
rect 6096 14116 6102 14118
rect 5794 14107 6102 14116
rect 36514 14172 36822 14181
rect 36514 14170 36520 14172
rect 36576 14170 36600 14172
rect 36656 14170 36680 14172
rect 36736 14170 36760 14172
rect 36816 14170 36822 14172
rect 36576 14118 36578 14170
rect 36758 14118 36760 14170
rect 36514 14116 36520 14118
rect 36576 14116 36600 14118
rect 36656 14116 36680 14118
rect 36736 14116 36760 14118
rect 36816 14116 36822 14118
rect 36514 14107 36822 14116
rect 67234 14172 67542 14181
rect 67234 14170 67240 14172
rect 67296 14170 67320 14172
rect 67376 14170 67400 14172
rect 67456 14170 67480 14172
rect 67536 14170 67542 14172
rect 67296 14118 67298 14170
rect 67478 14118 67480 14170
rect 67234 14116 67240 14118
rect 67296 14116 67320 14118
rect 67376 14116 67400 14118
rect 67456 14116 67480 14118
rect 67536 14116 67542 14118
rect 67234 14107 67542 14116
rect 5134 13628 5442 13637
rect 5134 13626 5140 13628
rect 5196 13626 5220 13628
rect 5276 13626 5300 13628
rect 5356 13626 5380 13628
rect 5436 13626 5442 13628
rect 5196 13574 5198 13626
rect 5378 13574 5380 13626
rect 5134 13572 5140 13574
rect 5196 13572 5220 13574
rect 5276 13572 5300 13574
rect 5356 13572 5380 13574
rect 5436 13572 5442 13574
rect 5134 13563 5442 13572
rect 35854 13628 36162 13637
rect 35854 13626 35860 13628
rect 35916 13626 35940 13628
rect 35996 13626 36020 13628
rect 36076 13626 36100 13628
rect 36156 13626 36162 13628
rect 35916 13574 35918 13626
rect 36098 13574 36100 13626
rect 35854 13572 35860 13574
rect 35916 13572 35940 13574
rect 35996 13572 36020 13574
rect 36076 13572 36100 13574
rect 36156 13572 36162 13574
rect 35854 13563 36162 13572
rect 66574 13628 66882 13637
rect 66574 13626 66580 13628
rect 66636 13626 66660 13628
rect 66716 13626 66740 13628
rect 66796 13626 66820 13628
rect 66876 13626 66882 13628
rect 66636 13574 66638 13626
rect 66818 13574 66820 13626
rect 66574 13572 66580 13574
rect 66636 13572 66660 13574
rect 66716 13572 66740 13574
rect 66796 13572 66820 13574
rect 66876 13572 66882 13574
rect 66574 13563 66882 13572
rect 5794 13084 6102 13093
rect 5794 13082 5800 13084
rect 5856 13082 5880 13084
rect 5936 13082 5960 13084
rect 6016 13082 6040 13084
rect 6096 13082 6102 13084
rect 5856 13030 5858 13082
rect 6038 13030 6040 13082
rect 5794 13028 5800 13030
rect 5856 13028 5880 13030
rect 5936 13028 5960 13030
rect 6016 13028 6040 13030
rect 6096 13028 6102 13030
rect 5794 13019 6102 13028
rect 36514 13084 36822 13093
rect 36514 13082 36520 13084
rect 36576 13082 36600 13084
rect 36656 13082 36680 13084
rect 36736 13082 36760 13084
rect 36816 13082 36822 13084
rect 36576 13030 36578 13082
rect 36758 13030 36760 13082
rect 36514 13028 36520 13030
rect 36576 13028 36600 13030
rect 36656 13028 36680 13030
rect 36736 13028 36760 13030
rect 36816 13028 36822 13030
rect 36514 13019 36822 13028
rect 67234 13084 67542 13093
rect 67234 13082 67240 13084
rect 67296 13082 67320 13084
rect 67376 13082 67400 13084
rect 67456 13082 67480 13084
rect 67536 13082 67542 13084
rect 67296 13030 67298 13082
rect 67478 13030 67480 13082
rect 67234 13028 67240 13030
rect 67296 13028 67320 13030
rect 67376 13028 67400 13030
rect 67456 13028 67480 13030
rect 67536 13028 67542 13030
rect 67234 13019 67542 13028
rect 5134 12540 5442 12549
rect 5134 12538 5140 12540
rect 5196 12538 5220 12540
rect 5276 12538 5300 12540
rect 5356 12538 5380 12540
rect 5436 12538 5442 12540
rect 5196 12486 5198 12538
rect 5378 12486 5380 12538
rect 5134 12484 5140 12486
rect 5196 12484 5220 12486
rect 5276 12484 5300 12486
rect 5356 12484 5380 12486
rect 5436 12484 5442 12486
rect 5134 12475 5442 12484
rect 35854 12540 36162 12549
rect 35854 12538 35860 12540
rect 35916 12538 35940 12540
rect 35996 12538 36020 12540
rect 36076 12538 36100 12540
rect 36156 12538 36162 12540
rect 35916 12486 35918 12538
rect 36098 12486 36100 12538
rect 35854 12484 35860 12486
rect 35916 12484 35940 12486
rect 35996 12484 36020 12486
rect 36076 12484 36100 12486
rect 36156 12484 36162 12486
rect 35854 12475 36162 12484
rect 66574 12540 66882 12549
rect 66574 12538 66580 12540
rect 66636 12538 66660 12540
rect 66716 12538 66740 12540
rect 66796 12538 66820 12540
rect 66876 12538 66882 12540
rect 66636 12486 66638 12538
rect 66818 12486 66820 12538
rect 66574 12484 66580 12486
rect 66636 12484 66660 12486
rect 66716 12484 66740 12486
rect 66796 12484 66820 12486
rect 66876 12484 66882 12486
rect 66574 12475 66882 12484
rect 5794 11996 6102 12005
rect 5794 11994 5800 11996
rect 5856 11994 5880 11996
rect 5936 11994 5960 11996
rect 6016 11994 6040 11996
rect 6096 11994 6102 11996
rect 5856 11942 5858 11994
rect 6038 11942 6040 11994
rect 5794 11940 5800 11942
rect 5856 11940 5880 11942
rect 5936 11940 5960 11942
rect 6016 11940 6040 11942
rect 6096 11940 6102 11942
rect 5794 11931 6102 11940
rect 36514 11996 36822 12005
rect 36514 11994 36520 11996
rect 36576 11994 36600 11996
rect 36656 11994 36680 11996
rect 36736 11994 36760 11996
rect 36816 11994 36822 11996
rect 36576 11942 36578 11994
rect 36758 11942 36760 11994
rect 36514 11940 36520 11942
rect 36576 11940 36600 11942
rect 36656 11940 36680 11942
rect 36736 11940 36760 11942
rect 36816 11940 36822 11942
rect 36514 11931 36822 11940
rect 67234 11996 67542 12005
rect 67234 11994 67240 11996
rect 67296 11994 67320 11996
rect 67376 11994 67400 11996
rect 67456 11994 67480 11996
rect 67536 11994 67542 11996
rect 67296 11942 67298 11994
rect 67478 11942 67480 11994
rect 67234 11940 67240 11942
rect 67296 11940 67320 11942
rect 67376 11940 67400 11942
rect 67456 11940 67480 11942
rect 67536 11940 67542 11942
rect 67234 11931 67542 11940
rect 5134 11452 5442 11461
rect 5134 11450 5140 11452
rect 5196 11450 5220 11452
rect 5276 11450 5300 11452
rect 5356 11450 5380 11452
rect 5436 11450 5442 11452
rect 5196 11398 5198 11450
rect 5378 11398 5380 11450
rect 5134 11396 5140 11398
rect 5196 11396 5220 11398
rect 5276 11396 5300 11398
rect 5356 11396 5380 11398
rect 5436 11396 5442 11398
rect 5134 11387 5442 11396
rect 35854 11452 36162 11461
rect 35854 11450 35860 11452
rect 35916 11450 35940 11452
rect 35996 11450 36020 11452
rect 36076 11450 36100 11452
rect 36156 11450 36162 11452
rect 35916 11398 35918 11450
rect 36098 11398 36100 11450
rect 35854 11396 35860 11398
rect 35916 11396 35940 11398
rect 35996 11396 36020 11398
rect 36076 11396 36100 11398
rect 36156 11396 36162 11398
rect 35854 11387 36162 11396
rect 66574 11452 66882 11461
rect 66574 11450 66580 11452
rect 66636 11450 66660 11452
rect 66716 11450 66740 11452
rect 66796 11450 66820 11452
rect 66876 11450 66882 11452
rect 66636 11398 66638 11450
rect 66818 11398 66820 11450
rect 66574 11396 66580 11398
rect 66636 11396 66660 11398
rect 66716 11396 66740 11398
rect 66796 11396 66820 11398
rect 66876 11396 66882 11398
rect 66574 11387 66882 11396
rect 5794 10908 6102 10917
rect 5794 10906 5800 10908
rect 5856 10906 5880 10908
rect 5936 10906 5960 10908
rect 6016 10906 6040 10908
rect 6096 10906 6102 10908
rect 5856 10854 5858 10906
rect 6038 10854 6040 10906
rect 5794 10852 5800 10854
rect 5856 10852 5880 10854
rect 5936 10852 5960 10854
rect 6016 10852 6040 10854
rect 6096 10852 6102 10854
rect 5794 10843 6102 10852
rect 36514 10908 36822 10917
rect 36514 10906 36520 10908
rect 36576 10906 36600 10908
rect 36656 10906 36680 10908
rect 36736 10906 36760 10908
rect 36816 10906 36822 10908
rect 36576 10854 36578 10906
rect 36758 10854 36760 10906
rect 36514 10852 36520 10854
rect 36576 10852 36600 10854
rect 36656 10852 36680 10854
rect 36736 10852 36760 10854
rect 36816 10852 36822 10854
rect 36514 10843 36822 10852
rect 67234 10908 67542 10917
rect 67234 10906 67240 10908
rect 67296 10906 67320 10908
rect 67376 10906 67400 10908
rect 67456 10906 67480 10908
rect 67536 10906 67542 10908
rect 67296 10854 67298 10906
rect 67478 10854 67480 10906
rect 67234 10852 67240 10854
rect 67296 10852 67320 10854
rect 67376 10852 67400 10854
rect 67456 10852 67480 10854
rect 67536 10852 67542 10854
rect 67234 10843 67542 10852
rect 5134 10364 5442 10373
rect 5134 10362 5140 10364
rect 5196 10362 5220 10364
rect 5276 10362 5300 10364
rect 5356 10362 5380 10364
rect 5436 10362 5442 10364
rect 5196 10310 5198 10362
rect 5378 10310 5380 10362
rect 5134 10308 5140 10310
rect 5196 10308 5220 10310
rect 5276 10308 5300 10310
rect 5356 10308 5380 10310
rect 5436 10308 5442 10310
rect 5134 10299 5442 10308
rect 35854 10364 36162 10373
rect 35854 10362 35860 10364
rect 35916 10362 35940 10364
rect 35996 10362 36020 10364
rect 36076 10362 36100 10364
rect 36156 10362 36162 10364
rect 35916 10310 35918 10362
rect 36098 10310 36100 10362
rect 35854 10308 35860 10310
rect 35916 10308 35940 10310
rect 35996 10308 36020 10310
rect 36076 10308 36100 10310
rect 36156 10308 36162 10310
rect 35854 10299 36162 10308
rect 66574 10364 66882 10373
rect 66574 10362 66580 10364
rect 66636 10362 66660 10364
rect 66716 10362 66740 10364
rect 66796 10362 66820 10364
rect 66876 10362 66882 10364
rect 66636 10310 66638 10362
rect 66818 10310 66820 10362
rect 66574 10308 66580 10310
rect 66636 10308 66660 10310
rect 66716 10308 66740 10310
rect 66796 10308 66820 10310
rect 66876 10308 66882 10310
rect 66574 10299 66882 10308
rect 5794 9820 6102 9829
rect 5794 9818 5800 9820
rect 5856 9818 5880 9820
rect 5936 9818 5960 9820
rect 6016 9818 6040 9820
rect 6096 9818 6102 9820
rect 5856 9766 5858 9818
rect 6038 9766 6040 9818
rect 5794 9764 5800 9766
rect 5856 9764 5880 9766
rect 5936 9764 5960 9766
rect 6016 9764 6040 9766
rect 6096 9764 6102 9766
rect 5794 9755 6102 9764
rect 36514 9820 36822 9829
rect 36514 9818 36520 9820
rect 36576 9818 36600 9820
rect 36656 9818 36680 9820
rect 36736 9818 36760 9820
rect 36816 9818 36822 9820
rect 36576 9766 36578 9818
rect 36758 9766 36760 9818
rect 36514 9764 36520 9766
rect 36576 9764 36600 9766
rect 36656 9764 36680 9766
rect 36736 9764 36760 9766
rect 36816 9764 36822 9766
rect 36514 9755 36822 9764
rect 67234 9820 67542 9829
rect 67234 9818 67240 9820
rect 67296 9818 67320 9820
rect 67376 9818 67400 9820
rect 67456 9818 67480 9820
rect 67536 9818 67542 9820
rect 67296 9766 67298 9818
rect 67478 9766 67480 9818
rect 67234 9764 67240 9766
rect 67296 9764 67320 9766
rect 67376 9764 67400 9766
rect 67456 9764 67480 9766
rect 67536 9764 67542 9766
rect 67234 9755 67542 9764
rect 5134 9276 5442 9285
rect 5134 9274 5140 9276
rect 5196 9274 5220 9276
rect 5276 9274 5300 9276
rect 5356 9274 5380 9276
rect 5436 9274 5442 9276
rect 5196 9222 5198 9274
rect 5378 9222 5380 9274
rect 5134 9220 5140 9222
rect 5196 9220 5220 9222
rect 5276 9220 5300 9222
rect 5356 9220 5380 9222
rect 5436 9220 5442 9222
rect 5134 9211 5442 9220
rect 35854 9276 36162 9285
rect 35854 9274 35860 9276
rect 35916 9274 35940 9276
rect 35996 9274 36020 9276
rect 36076 9274 36100 9276
rect 36156 9274 36162 9276
rect 35916 9222 35918 9274
rect 36098 9222 36100 9274
rect 35854 9220 35860 9222
rect 35916 9220 35940 9222
rect 35996 9220 36020 9222
rect 36076 9220 36100 9222
rect 36156 9220 36162 9222
rect 35854 9211 36162 9220
rect 66574 9276 66882 9285
rect 66574 9274 66580 9276
rect 66636 9274 66660 9276
rect 66716 9274 66740 9276
rect 66796 9274 66820 9276
rect 66876 9274 66882 9276
rect 66636 9222 66638 9274
rect 66818 9222 66820 9274
rect 66574 9220 66580 9222
rect 66636 9220 66660 9222
rect 66716 9220 66740 9222
rect 66796 9220 66820 9222
rect 66876 9220 66882 9222
rect 66574 9211 66882 9220
rect 5794 8732 6102 8741
rect 5794 8730 5800 8732
rect 5856 8730 5880 8732
rect 5936 8730 5960 8732
rect 6016 8730 6040 8732
rect 6096 8730 6102 8732
rect 5856 8678 5858 8730
rect 6038 8678 6040 8730
rect 5794 8676 5800 8678
rect 5856 8676 5880 8678
rect 5936 8676 5960 8678
rect 6016 8676 6040 8678
rect 6096 8676 6102 8678
rect 5794 8667 6102 8676
rect 36514 8732 36822 8741
rect 36514 8730 36520 8732
rect 36576 8730 36600 8732
rect 36656 8730 36680 8732
rect 36736 8730 36760 8732
rect 36816 8730 36822 8732
rect 36576 8678 36578 8730
rect 36758 8678 36760 8730
rect 36514 8676 36520 8678
rect 36576 8676 36600 8678
rect 36656 8676 36680 8678
rect 36736 8676 36760 8678
rect 36816 8676 36822 8678
rect 36514 8667 36822 8676
rect 67234 8732 67542 8741
rect 67234 8730 67240 8732
rect 67296 8730 67320 8732
rect 67376 8730 67400 8732
rect 67456 8730 67480 8732
rect 67536 8730 67542 8732
rect 67296 8678 67298 8730
rect 67478 8678 67480 8730
rect 67234 8676 67240 8678
rect 67296 8676 67320 8678
rect 67376 8676 67400 8678
rect 67456 8676 67480 8678
rect 67536 8676 67542 8678
rect 67234 8667 67542 8676
rect 5134 8188 5442 8197
rect 5134 8186 5140 8188
rect 5196 8186 5220 8188
rect 5276 8186 5300 8188
rect 5356 8186 5380 8188
rect 5436 8186 5442 8188
rect 5196 8134 5198 8186
rect 5378 8134 5380 8186
rect 5134 8132 5140 8134
rect 5196 8132 5220 8134
rect 5276 8132 5300 8134
rect 5356 8132 5380 8134
rect 5436 8132 5442 8134
rect 5134 8123 5442 8132
rect 35854 8188 36162 8197
rect 35854 8186 35860 8188
rect 35916 8186 35940 8188
rect 35996 8186 36020 8188
rect 36076 8186 36100 8188
rect 36156 8186 36162 8188
rect 35916 8134 35918 8186
rect 36098 8134 36100 8186
rect 35854 8132 35860 8134
rect 35916 8132 35940 8134
rect 35996 8132 36020 8134
rect 36076 8132 36100 8134
rect 36156 8132 36162 8134
rect 35854 8123 36162 8132
rect 66574 8188 66882 8197
rect 66574 8186 66580 8188
rect 66636 8186 66660 8188
rect 66716 8186 66740 8188
rect 66796 8186 66820 8188
rect 66876 8186 66882 8188
rect 66636 8134 66638 8186
rect 66818 8134 66820 8186
rect 66574 8132 66580 8134
rect 66636 8132 66660 8134
rect 66716 8132 66740 8134
rect 66796 8132 66820 8134
rect 66876 8132 66882 8134
rect 66574 8123 66882 8132
rect 5794 7644 6102 7653
rect 5794 7642 5800 7644
rect 5856 7642 5880 7644
rect 5936 7642 5960 7644
rect 6016 7642 6040 7644
rect 6096 7642 6102 7644
rect 5856 7590 5858 7642
rect 6038 7590 6040 7642
rect 5794 7588 5800 7590
rect 5856 7588 5880 7590
rect 5936 7588 5960 7590
rect 6016 7588 6040 7590
rect 6096 7588 6102 7590
rect 5794 7579 6102 7588
rect 36514 7644 36822 7653
rect 36514 7642 36520 7644
rect 36576 7642 36600 7644
rect 36656 7642 36680 7644
rect 36736 7642 36760 7644
rect 36816 7642 36822 7644
rect 36576 7590 36578 7642
rect 36758 7590 36760 7642
rect 36514 7588 36520 7590
rect 36576 7588 36600 7590
rect 36656 7588 36680 7590
rect 36736 7588 36760 7590
rect 36816 7588 36822 7590
rect 36514 7579 36822 7588
rect 67234 7644 67542 7653
rect 67234 7642 67240 7644
rect 67296 7642 67320 7644
rect 67376 7642 67400 7644
rect 67456 7642 67480 7644
rect 67536 7642 67542 7644
rect 67296 7590 67298 7642
rect 67478 7590 67480 7642
rect 67234 7588 67240 7590
rect 67296 7588 67320 7590
rect 67376 7588 67400 7590
rect 67456 7588 67480 7590
rect 67536 7588 67542 7590
rect 67234 7579 67542 7588
rect 5134 7100 5442 7109
rect 5134 7098 5140 7100
rect 5196 7098 5220 7100
rect 5276 7098 5300 7100
rect 5356 7098 5380 7100
rect 5436 7098 5442 7100
rect 5196 7046 5198 7098
rect 5378 7046 5380 7098
rect 5134 7044 5140 7046
rect 5196 7044 5220 7046
rect 5276 7044 5300 7046
rect 5356 7044 5380 7046
rect 5436 7044 5442 7046
rect 5134 7035 5442 7044
rect 35854 7100 36162 7109
rect 35854 7098 35860 7100
rect 35916 7098 35940 7100
rect 35996 7098 36020 7100
rect 36076 7098 36100 7100
rect 36156 7098 36162 7100
rect 35916 7046 35918 7098
rect 36098 7046 36100 7098
rect 35854 7044 35860 7046
rect 35916 7044 35940 7046
rect 35996 7044 36020 7046
rect 36076 7044 36100 7046
rect 36156 7044 36162 7046
rect 35854 7035 36162 7044
rect 66574 7100 66882 7109
rect 66574 7098 66580 7100
rect 66636 7098 66660 7100
rect 66716 7098 66740 7100
rect 66796 7098 66820 7100
rect 66876 7098 66882 7100
rect 66636 7046 66638 7098
rect 66818 7046 66820 7098
rect 66574 7044 66580 7046
rect 66636 7044 66660 7046
rect 66716 7044 66740 7046
rect 66796 7044 66820 7046
rect 66876 7044 66882 7046
rect 66574 7035 66882 7044
rect 5794 6556 6102 6565
rect 5794 6554 5800 6556
rect 5856 6554 5880 6556
rect 5936 6554 5960 6556
rect 6016 6554 6040 6556
rect 6096 6554 6102 6556
rect 5856 6502 5858 6554
rect 6038 6502 6040 6554
rect 5794 6500 5800 6502
rect 5856 6500 5880 6502
rect 5936 6500 5960 6502
rect 6016 6500 6040 6502
rect 6096 6500 6102 6502
rect 5794 6491 6102 6500
rect 36514 6556 36822 6565
rect 36514 6554 36520 6556
rect 36576 6554 36600 6556
rect 36656 6554 36680 6556
rect 36736 6554 36760 6556
rect 36816 6554 36822 6556
rect 36576 6502 36578 6554
rect 36758 6502 36760 6554
rect 36514 6500 36520 6502
rect 36576 6500 36600 6502
rect 36656 6500 36680 6502
rect 36736 6500 36760 6502
rect 36816 6500 36822 6502
rect 36514 6491 36822 6500
rect 67234 6556 67542 6565
rect 67234 6554 67240 6556
rect 67296 6554 67320 6556
rect 67376 6554 67400 6556
rect 67456 6554 67480 6556
rect 67536 6554 67542 6556
rect 67296 6502 67298 6554
rect 67478 6502 67480 6554
rect 67234 6500 67240 6502
rect 67296 6500 67320 6502
rect 67376 6500 67400 6502
rect 67456 6500 67480 6502
rect 67536 6500 67542 6502
rect 67234 6491 67542 6500
rect 5134 6012 5442 6021
rect 5134 6010 5140 6012
rect 5196 6010 5220 6012
rect 5276 6010 5300 6012
rect 5356 6010 5380 6012
rect 5436 6010 5442 6012
rect 5196 5958 5198 6010
rect 5378 5958 5380 6010
rect 5134 5956 5140 5958
rect 5196 5956 5220 5958
rect 5276 5956 5300 5958
rect 5356 5956 5380 5958
rect 5436 5956 5442 5958
rect 5134 5947 5442 5956
rect 35854 6012 36162 6021
rect 35854 6010 35860 6012
rect 35916 6010 35940 6012
rect 35996 6010 36020 6012
rect 36076 6010 36100 6012
rect 36156 6010 36162 6012
rect 35916 5958 35918 6010
rect 36098 5958 36100 6010
rect 35854 5956 35860 5958
rect 35916 5956 35940 5958
rect 35996 5956 36020 5958
rect 36076 5956 36100 5958
rect 36156 5956 36162 5958
rect 35854 5947 36162 5956
rect 66574 6012 66882 6021
rect 66574 6010 66580 6012
rect 66636 6010 66660 6012
rect 66716 6010 66740 6012
rect 66796 6010 66820 6012
rect 66876 6010 66882 6012
rect 66636 5958 66638 6010
rect 66818 5958 66820 6010
rect 66574 5956 66580 5958
rect 66636 5956 66660 5958
rect 66716 5956 66740 5958
rect 66796 5956 66820 5958
rect 66876 5956 66882 5958
rect 66574 5947 66882 5956
rect 5794 5468 6102 5477
rect 5794 5466 5800 5468
rect 5856 5466 5880 5468
rect 5936 5466 5960 5468
rect 6016 5466 6040 5468
rect 6096 5466 6102 5468
rect 5856 5414 5858 5466
rect 6038 5414 6040 5466
rect 5794 5412 5800 5414
rect 5856 5412 5880 5414
rect 5936 5412 5960 5414
rect 6016 5412 6040 5414
rect 6096 5412 6102 5414
rect 5794 5403 6102 5412
rect 36514 5468 36822 5477
rect 36514 5466 36520 5468
rect 36576 5466 36600 5468
rect 36656 5466 36680 5468
rect 36736 5466 36760 5468
rect 36816 5466 36822 5468
rect 36576 5414 36578 5466
rect 36758 5414 36760 5466
rect 36514 5412 36520 5414
rect 36576 5412 36600 5414
rect 36656 5412 36680 5414
rect 36736 5412 36760 5414
rect 36816 5412 36822 5414
rect 36514 5403 36822 5412
rect 67234 5468 67542 5477
rect 67234 5466 67240 5468
rect 67296 5466 67320 5468
rect 67376 5466 67400 5468
rect 67456 5466 67480 5468
rect 67536 5466 67542 5468
rect 67296 5414 67298 5466
rect 67478 5414 67480 5466
rect 67234 5412 67240 5414
rect 67296 5412 67320 5414
rect 67376 5412 67400 5414
rect 67456 5412 67480 5414
rect 67536 5412 67542 5414
rect 67234 5403 67542 5412
rect 5134 4924 5442 4933
rect 5134 4922 5140 4924
rect 5196 4922 5220 4924
rect 5276 4922 5300 4924
rect 5356 4922 5380 4924
rect 5436 4922 5442 4924
rect 5196 4870 5198 4922
rect 5378 4870 5380 4922
rect 5134 4868 5140 4870
rect 5196 4868 5220 4870
rect 5276 4868 5300 4870
rect 5356 4868 5380 4870
rect 5436 4868 5442 4870
rect 5134 4859 5442 4868
rect 35854 4924 36162 4933
rect 35854 4922 35860 4924
rect 35916 4922 35940 4924
rect 35996 4922 36020 4924
rect 36076 4922 36100 4924
rect 36156 4922 36162 4924
rect 35916 4870 35918 4922
rect 36098 4870 36100 4922
rect 35854 4868 35860 4870
rect 35916 4868 35940 4870
rect 35996 4868 36020 4870
rect 36076 4868 36100 4870
rect 36156 4868 36162 4870
rect 35854 4859 36162 4868
rect 66574 4924 66882 4933
rect 66574 4922 66580 4924
rect 66636 4922 66660 4924
rect 66716 4922 66740 4924
rect 66796 4922 66820 4924
rect 66876 4922 66882 4924
rect 66636 4870 66638 4922
rect 66818 4870 66820 4922
rect 66574 4868 66580 4870
rect 66636 4868 66660 4870
rect 66716 4868 66740 4870
rect 66796 4868 66820 4870
rect 66876 4868 66882 4870
rect 66574 4859 66882 4868
rect 5794 4380 6102 4389
rect 5794 4378 5800 4380
rect 5856 4378 5880 4380
rect 5936 4378 5960 4380
rect 6016 4378 6040 4380
rect 6096 4378 6102 4380
rect 5856 4326 5858 4378
rect 6038 4326 6040 4378
rect 5794 4324 5800 4326
rect 5856 4324 5880 4326
rect 5936 4324 5960 4326
rect 6016 4324 6040 4326
rect 6096 4324 6102 4326
rect 5794 4315 6102 4324
rect 36514 4380 36822 4389
rect 36514 4378 36520 4380
rect 36576 4378 36600 4380
rect 36656 4378 36680 4380
rect 36736 4378 36760 4380
rect 36816 4378 36822 4380
rect 36576 4326 36578 4378
rect 36758 4326 36760 4378
rect 36514 4324 36520 4326
rect 36576 4324 36600 4326
rect 36656 4324 36680 4326
rect 36736 4324 36760 4326
rect 36816 4324 36822 4326
rect 36514 4315 36822 4324
rect 67234 4380 67542 4389
rect 67234 4378 67240 4380
rect 67296 4378 67320 4380
rect 67376 4378 67400 4380
rect 67456 4378 67480 4380
rect 67536 4378 67542 4380
rect 67296 4326 67298 4378
rect 67478 4326 67480 4378
rect 67234 4324 67240 4326
rect 67296 4324 67320 4326
rect 67376 4324 67400 4326
rect 67456 4324 67480 4326
rect 67536 4324 67542 4326
rect 67234 4315 67542 4324
rect 5134 3836 5442 3845
rect 5134 3834 5140 3836
rect 5196 3834 5220 3836
rect 5276 3834 5300 3836
rect 5356 3834 5380 3836
rect 5436 3834 5442 3836
rect 5196 3782 5198 3834
rect 5378 3782 5380 3834
rect 5134 3780 5140 3782
rect 5196 3780 5220 3782
rect 5276 3780 5300 3782
rect 5356 3780 5380 3782
rect 5436 3780 5442 3782
rect 5134 3771 5442 3780
rect 35854 3836 36162 3845
rect 35854 3834 35860 3836
rect 35916 3834 35940 3836
rect 35996 3834 36020 3836
rect 36076 3834 36100 3836
rect 36156 3834 36162 3836
rect 35916 3782 35918 3834
rect 36098 3782 36100 3834
rect 35854 3780 35860 3782
rect 35916 3780 35940 3782
rect 35996 3780 36020 3782
rect 36076 3780 36100 3782
rect 36156 3780 36162 3782
rect 35854 3771 36162 3780
rect 66574 3836 66882 3845
rect 66574 3834 66580 3836
rect 66636 3834 66660 3836
rect 66716 3834 66740 3836
rect 66796 3834 66820 3836
rect 66876 3834 66882 3836
rect 66636 3782 66638 3834
rect 66818 3782 66820 3834
rect 66574 3780 66580 3782
rect 66636 3780 66660 3782
rect 66716 3780 66740 3782
rect 66796 3780 66820 3782
rect 66876 3780 66882 3782
rect 66574 3771 66882 3780
rect 5794 3292 6102 3301
rect 5794 3290 5800 3292
rect 5856 3290 5880 3292
rect 5936 3290 5960 3292
rect 6016 3290 6040 3292
rect 6096 3290 6102 3292
rect 5856 3238 5858 3290
rect 6038 3238 6040 3290
rect 5794 3236 5800 3238
rect 5856 3236 5880 3238
rect 5936 3236 5960 3238
rect 6016 3236 6040 3238
rect 6096 3236 6102 3238
rect 5794 3227 6102 3236
rect 36514 3292 36822 3301
rect 36514 3290 36520 3292
rect 36576 3290 36600 3292
rect 36656 3290 36680 3292
rect 36736 3290 36760 3292
rect 36816 3290 36822 3292
rect 36576 3238 36578 3290
rect 36758 3238 36760 3290
rect 36514 3236 36520 3238
rect 36576 3236 36600 3238
rect 36656 3236 36680 3238
rect 36736 3236 36760 3238
rect 36816 3236 36822 3238
rect 36514 3227 36822 3236
rect 67234 3292 67542 3301
rect 67234 3290 67240 3292
rect 67296 3290 67320 3292
rect 67376 3290 67400 3292
rect 67456 3290 67480 3292
rect 67536 3290 67542 3292
rect 67296 3238 67298 3290
rect 67478 3238 67480 3290
rect 67234 3236 67240 3238
rect 67296 3236 67320 3238
rect 67376 3236 67400 3238
rect 67456 3236 67480 3238
rect 67536 3236 67542 3238
rect 67234 3227 67542 3236
rect 5134 2748 5442 2757
rect 5134 2746 5140 2748
rect 5196 2746 5220 2748
rect 5276 2746 5300 2748
rect 5356 2746 5380 2748
rect 5436 2746 5442 2748
rect 5196 2694 5198 2746
rect 5378 2694 5380 2746
rect 5134 2692 5140 2694
rect 5196 2692 5220 2694
rect 5276 2692 5300 2694
rect 5356 2692 5380 2694
rect 5436 2692 5442 2694
rect 5134 2683 5442 2692
rect 35854 2748 36162 2757
rect 35854 2746 35860 2748
rect 35916 2746 35940 2748
rect 35996 2746 36020 2748
rect 36076 2746 36100 2748
rect 36156 2746 36162 2748
rect 35916 2694 35918 2746
rect 36098 2694 36100 2746
rect 35854 2692 35860 2694
rect 35916 2692 35940 2694
rect 35996 2692 36020 2694
rect 36076 2692 36100 2694
rect 36156 2692 36162 2694
rect 35854 2683 36162 2692
rect 66574 2748 66882 2757
rect 66574 2746 66580 2748
rect 66636 2746 66660 2748
rect 66716 2746 66740 2748
rect 66796 2746 66820 2748
rect 66876 2746 66882 2748
rect 66636 2694 66638 2746
rect 66818 2694 66820 2746
rect 66574 2692 66580 2694
rect 66636 2692 66660 2694
rect 66716 2692 66740 2694
rect 66796 2692 66820 2694
rect 66876 2692 66882 2694
rect 66574 2683 66882 2692
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 41880 2440 41932 2446
rect 41880 2382 41932 2388
rect 42524 2440 42576 2446
rect 42524 2382 42576 2388
rect 44456 2440 44508 2446
rect 44456 2382 44508 2388
rect 52184 2440 52236 2446
rect 52184 2382 52236 2388
rect 57980 2440 58032 2446
rect 57980 2382 58032 2388
rect 59268 2440 59320 2446
rect 59268 2382 59320 2388
rect 5794 2204 6102 2213
rect 5794 2202 5800 2204
rect 5856 2202 5880 2204
rect 5936 2202 5960 2204
rect 6016 2202 6040 2204
rect 6096 2202 6102 2204
rect 5856 2150 5858 2202
rect 6038 2150 6040 2202
rect 5794 2148 5800 2150
rect 5856 2148 5880 2150
rect 5936 2148 5960 2150
rect 6016 2148 6040 2150
rect 6096 2148 6102 2150
rect 5794 2139 6102 2148
rect 22572 800 22600 2382
rect 23216 800 23244 2382
rect 33520 800 33548 2382
rect 36514 2204 36822 2213
rect 36514 2202 36520 2204
rect 36576 2202 36600 2204
rect 36656 2202 36680 2204
rect 36736 2202 36760 2204
rect 36816 2202 36822 2204
rect 36576 2150 36578 2202
rect 36758 2150 36760 2202
rect 36514 2148 36520 2150
rect 36576 2148 36600 2150
rect 36656 2148 36680 2150
rect 36736 2148 36760 2150
rect 36816 2148 36822 2150
rect 36514 2139 36822 2148
rect 41892 800 41920 2382
rect 42536 800 42564 2382
rect 44468 800 44496 2382
rect 52196 800 52224 2382
rect 57992 800 58020 2382
rect 59280 800 59308 2382
rect 67234 2204 67542 2213
rect 67234 2202 67240 2204
rect 67296 2202 67320 2204
rect 67376 2202 67400 2204
rect 67456 2202 67480 2204
rect 67536 2202 67542 2204
rect 67296 2150 67298 2202
rect 67478 2150 67480 2202
rect 67234 2148 67240 2150
rect 67296 2148 67320 2150
rect 67376 2148 67400 2150
rect 67456 2148 67480 2150
rect 67536 2148 67542 2150
rect 67234 2139 67542 2148
rect 18 0 74 800
rect 662 0 718 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 33506 0 33562 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 44454 0 44510 800
rect 52182 0 52238 800
rect 57978 0 58034 800
rect 59266 0 59322 800
<< via2 >>
rect 5140 77818 5196 77820
rect 5220 77818 5276 77820
rect 5300 77818 5356 77820
rect 5380 77818 5436 77820
rect 5140 77766 5186 77818
rect 5186 77766 5196 77818
rect 5220 77766 5250 77818
rect 5250 77766 5262 77818
rect 5262 77766 5276 77818
rect 5300 77766 5314 77818
rect 5314 77766 5326 77818
rect 5326 77766 5356 77818
rect 5380 77766 5390 77818
rect 5390 77766 5436 77818
rect 5140 77764 5196 77766
rect 5220 77764 5276 77766
rect 5300 77764 5356 77766
rect 5380 77764 5436 77766
rect 35860 77818 35916 77820
rect 35940 77818 35996 77820
rect 36020 77818 36076 77820
rect 36100 77818 36156 77820
rect 35860 77766 35906 77818
rect 35906 77766 35916 77818
rect 35940 77766 35970 77818
rect 35970 77766 35982 77818
rect 35982 77766 35996 77818
rect 36020 77766 36034 77818
rect 36034 77766 36046 77818
rect 36046 77766 36076 77818
rect 36100 77766 36110 77818
rect 36110 77766 36156 77818
rect 35860 77764 35916 77766
rect 35940 77764 35996 77766
rect 36020 77764 36076 77766
rect 36100 77764 36156 77766
rect 66580 77818 66636 77820
rect 66660 77818 66716 77820
rect 66740 77818 66796 77820
rect 66820 77818 66876 77820
rect 66580 77766 66626 77818
rect 66626 77766 66636 77818
rect 66660 77766 66690 77818
rect 66690 77766 66702 77818
rect 66702 77766 66716 77818
rect 66740 77766 66754 77818
rect 66754 77766 66766 77818
rect 66766 77766 66796 77818
rect 66820 77766 66830 77818
rect 66830 77766 66876 77818
rect 66580 77764 66636 77766
rect 66660 77764 66716 77766
rect 66740 77764 66796 77766
rect 66820 77764 66876 77766
rect 5800 77274 5856 77276
rect 5880 77274 5936 77276
rect 5960 77274 6016 77276
rect 6040 77274 6096 77276
rect 5800 77222 5846 77274
rect 5846 77222 5856 77274
rect 5880 77222 5910 77274
rect 5910 77222 5922 77274
rect 5922 77222 5936 77274
rect 5960 77222 5974 77274
rect 5974 77222 5986 77274
rect 5986 77222 6016 77274
rect 6040 77222 6050 77274
rect 6050 77222 6096 77274
rect 5800 77220 5856 77222
rect 5880 77220 5936 77222
rect 5960 77220 6016 77222
rect 6040 77220 6096 77222
rect 36520 77274 36576 77276
rect 36600 77274 36656 77276
rect 36680 77274 36736 77276
rect 36760 77274 36816 77276
rect 36520 77222 36566 77274
rect 36566 77222 36576 77274
rect 36600 77222 36630 77274
rect 36630 77222 36642 77274
rect 36642 77222 36656 77274
rect 36680 77222 36694 77274
rect 36694 77222 36706 77274
rect 36706 77222 36736 77274
rect 36760 77222 36770 77274
rect 36770 77222 36816 77274
rect 36520 77220 36576 77222
rect 36600 77220 36656 77222
rect 36680 77220 36736 77222
rect 36760 77220 36816 77222
rect 67240 77274 67296 77276
rect 67320 77274 67376 77276
rect 67400 77274 67456 77276
rect 67480 77274 67536 77276
rect 67240 77222 67286 77274
rect 67286 77222 67296 77274
rect 67320 77222 67350 77274
rect 67350 77222 67362 77274
rect 67362 77222 67376 77274
rect 67400 77222 67414 77274
rect 67414 77222 67426 77274
rect 67426 77222 67456 77274
rect 67480 77222 67490 77274
rect 67490 77222 67536 77274
rect 67240 77220 67296 77222
rect 67320 77220 67376 77222
rect 67400 77220 67456 77222
rect 67480 77220 67536 77222
rect 5140 76730 5196 76732
rect 5220 76730 5276 76732
rect 5300 76730 5356 76732
rect 5380 76730 5436 76732
rect 5140 76678 5186 76730
rect 5186 76678 5196 76730
rect 5220 76678 5250 76730
rect 5250 76678 5262 76730
rect 5262 76678 5276 76730
rect 5300 76678 5314 76730
rect 5314 76678 5326 76730
rect 5326 76678 5356 76730
rect 5380 76678 5390 76730
rect 5390 76678 5436 76730
rect 5140 76676 5196 76678
rect 5220 76676 5276 76678
rect 5300 76676 5356 76678
rect 5380 76676 5436 76678
rect 35860 76730 35916 76732
rect 35940 76730 35996 76732
rect 36020 76730 36076 76732
rect 36100 76730 36156 76732
rect 35860 76678 35906 76730
rect 35906 76678 35916 76730
rect 35940 76678 35970 76730
rect 35970 76678 35982 76730
rect 35982 76678 35996 76730
rect 36020 76678 36034 76730
rect 36034 76678 36046 76730
rect 36046 76678 36076 76730
rect 36100 76678 36110 76730
rect 36110 76678 36156 76730
rect 35860 76676 35916 76678
rect 35940 76676 35996 76678
rect 36020 76676 36076 76678
rect 36100 76676 36156 76678
rect 66580 76730 66636 76732
rect 66660 76730 66716 76732
rect 66740 76730 66796 76732
rect 66820 76730 66876 76732
rect 66580 76678 66626 76730
rect 66626 76678 66636 76730
rect 66660 76678 66690 76730
rect 66690 76678 66702 76730
rect 66702 76678 66716 76730
rect 66740 76678 66754 76730
rect 66754 76678 66766 76730
rect 66766 76678 66796 76730
rect 66820 76678 66830 76730
rect 66830 76678 66876 76730
rect 66580 76676 66636 76678
rect 66660 76676 66716 76678
rect 66740 76676 66796 76678
rect 66820 76676 66876 76678
rect 5800 76186 5856 76188
rect 5880 76186 5936 76188
rect 5960 76186 6016 76188
rect 6040 76186 6096 76188
rect 5800 76134 5846 76186
rect 5846 76134 5856 76186
rect 5880 76134 5910 76186
rect 5910 76134 5922 76186
rect 5922 76134 5936 76186
rect 5960 76134 5974 76186
rect 5974 76134 5986 76186
rect 5986 76134 6016 76186
rect 6040 76134 6050 76186
rect 6050 76134 6096 76186
rect 5800 76132 5856 76134
rect 5880 76132 5936 76134
rect 5960 76132 6016 76134
rect 6040 76132 6096 76134
rect 36520 76186 36576 76188
rect 36600 76186 36656 76188
rect 36680 76186 36736 76188
rect 36760 76186 36816 76188
rect 36520 76134 36566 76186
rect 36566 76134 36576 76186
rect 36600 76134 36630 76186
rect 36630 76134 36642 76186
rect 36642 76134 36656 76186
rect 36680 76134 36694 76186
rect 36694 76134 36706 76186
rect 36706 76134 36736 76186
rect 36760 76134 36770 76186
rect 36770 76134 36816 76186
rect 36520 76132 36576 76134
rect 36600 76132 36656 76134
rect 36680 76132 36736 76134
rect 36760 76132 36816 76134
rect 67240 76186 67296 76188
rect 67320 76186 67376 76188
rect 67400 76186 67456 76188
rect 67480 76186 67536 76188
rect 67240 76134 67286 76186
rect 67286 76134 67296 76186
rect 67320 76134 67350 76186
rect 67350 76134 67362 76186
rect 67362 76134 67376 76186
rect 67400 76134 67414 76186
rect 67414 76134 67426 76186
rect 67426 76134 67456 76186
rect 67480 76134 67490 76186
rect 67490 76134 67536 76186
rect 67240 76132 67296 76134
rect 67320 76132 67376 76134
rect 67400 76132 67456 76134
rect 67480 76132 67536 76134
rect 5140 75642 5196 75644
rect 5220 75642 5276 75644
rect 5300 75642 5356 75644
rect 5380 75642 5436 75644
rect 5140 75590 5186 75642
rect 5186 75590 5196 75642
rect 5220 75590 5250 75642
rect 5250 75590 5262 75642
rect 5262 75590 5276 75642
rect 5300 75590 5314 75642
rect 5314 75590 5326 75642
rect 5326 75590 5356 75642
rect 5380 75590 5390 75642
rect 5390 75590 5436 75642
rect 5140 75588 5196 75590
rect 5220 75588 5276 75590
rect 5300 75588 5356 75590
rect 5380 75588 5436 75590
rect 35860 75642 35916 75644
rect 35940 75642 35996 75644
rect 36020 75642 36076 75644
rect 36100 75642 36156 75644
rect 35860 75590 35906 75642
rect 35906 75590 35916 75642
rect 35940 75590 35970 75642
rect 35970 75590 35982 75642
rect 35982 75590 35996 75642
rect 36020 75590 36034 75642
rect 36034 75590 36046 75642
rect 36046 75590 36076 75642
rect 36100 75590 36110 75642
rect 36110 75590 36156 75642
rect 35860 75588 35916 75590
rect 35940 75588 35996 75590
rect 36020 75588 36076 75590
rect 36100 75588 36156 75590
rect 66580 75642 66636 75644
rect 66660 75642 66716 75644
rect 66740 75642 66796 75644
rect 66820 75642 66876 75644
rect 66580 75590 66626 75642
rect 66626 75590 66636 75642
rect 66660 75590 66690 75642
rect 66690 75590 66702 75642
rect 66702 75590 66716 75642
rect 66740 75590 66754 75642
rect 66754 75590 66766 75642
rect 66766 75590 66796 75642
rect 66820 75590 66830 75642
rect 66830 75590 66876 75642
rect 66580 75588 66636 75590
rect 66660 75588 66716 75590
rect 66740 75588 66796 75590
rect 66820 75588 66876 75590
rect 5800 75098 5856 75100
rect 5880 75098 5936 75100
rect 5960 75098 6016 75100
rect 6040 75098 6096 75100
rect 5800 75046 5846 75098
rect 5846 75046 5856 75098
rect 5880 75046 5910 75098
rect 5910 75046 5922 75098
rect 5922 75046 5936 75098
rect 5960 75046 5974 75098
rect 5974 75046 5986 75098
rect 5986 75046 6016 75098
rect 6040 75046 6050 75098
rect 6050 75046 6096 75098
rect 5800 75044 5856 75046
rect 5880 75044 5936 75046
rect 5960 75044 6016 75046
rect 6040 75044 6096 75046
rect 36520 75098 36576 75100
rect 36600 75098 36656 75100
rect 36680 75098 36736 75100
rect 36760 75098 36816 75100
rect 36520 75046 36566 75098
rect 36566 75046 36576 75098
rect 36600 75046 36630 75098
rect 36630 75046 36642 75098
rect 36642 75046 36656 75098
rect 36680 75046 36694 75098
rect 36694 75046 36706 75098
rect 36706 75046 36736 75098
rect 36760 75046 36770 75098
rect 36770 75046 36816 75098
rect 36520 75044 36576 75046
rect 36600 75044 36656 75046
rect 36680 75044 36736 75046
rect 36760 75044 36816 75046
rect 67240 75098 67296 75100
rect 67320 75098 67376 75100
rect 67400 75098 67456 75100
rect 67480 75098 67536 75100
rect 67240 75046 67286 75098
rect 67286 75046 67296 75098
rect 67320 75046 67350 75098
rect 67350 75046 67362 75098
rect 67362 75046 67376 75098
rect 67400 75046 67414 75098
rect 67414 75046 67426 75098
rect 67426 75046 67456 75098
rect 67480 75046 67490 75098
rect 67490 75046 67536 75098
rect 67240 75044 67296 75046
rect 67320 75044 67376 75046
rect 67400 75044 67456 75046
rect 67480 75044 67536 75046
rect 5140 74554 5196 74556
rect 5220 74554 5276 74556
rect 5300 74554 5356 74556
rect 5380 74554 5436 74556
rect 5140 74502 5186 74554
rect 5186 74502 5196 74554
rect 5220 74502 5250 74554
rect 5250 74502 5262 74554
rect 5262 74502 5276 74554
rect 5300 74502 5314 74554
rect 5314 74502 5326 74554
rect 5326 74502 5356 74554
rect 5380 74502 5390 74554
rect 5390 74502 5436 74554
rect 5140 74500 5196 74502
rect 5220 74500 5276 74502
rect 5300 74500 5356 74502
rect 5380 74500 5436 74502
rect 35860 74554 35916 74556
rect 35940 74554 35996 74556
rect 36020 74554 36076 74556
rect 36100 74554 36156 74556
rect 35860 74502 35906 74554
rect 35906 74502 35916 74554
rect 35940 74502 35970 74554
rect 35970 74502 35982 74554
rect 35982 74502 35996 74554
rect 36020 74502 36034 74554
rect 36034 74502 36046 74554
rect 36046 74502 36076 74554
rect 36100 74502 36110 74554
rect 36110 74502 36156 74554
rect 35860 74500 35916 74502
rect 35940 74500 35996 74502
rect 36020 74500 36076 74502
rect 36100 74500 36156 74502
rect 66580 74554 66636 74556
rect 66660 74554 66716 74556
rect 66740 74554 66796 74556
rect 66820 74554 66876 74556
rect 66580 74502 66626 74554
rect 66626 74502 66636 74554
rect 66660 74502 66690 74554
rect 66690 74502 66702 74554
rect 66702 74502 66716 74554
rect 66740 74502 66754 74554
rect 66754 74502 66766 74554
rect 66766 74502 66796 74554
rect 66820 74502 66830 74554
rect 66830 74502 66876 74554
rect 66580 74500 66636 74502
rect 66660 74500 66716 74502
rect 66740 74500 66796 74502
rect 66820 74500 66876 74502
rect 5800 74010 5856 74012
rect 5880 74010 5936 74012
rect 5960 74010 6016 74012
rect 6040 74010 6096 74012
rect 5800 73958 5846 74010
rect 5846 73958 5856 74010
rect 5880 73958 5910 74010
rect 5910 73958 5922 74010
rect 5922 73958 5936 74010
rect 5960 73958 5974 74010
rect 5974 73958 5986 74010
rect 5986 73958 6016 74010
rect 6040 73958 6050 74010
rect 6050 73958 6096 74010
rect 5800 73956 5856 73958
rect 5880 73956 5936 73958
rect 5960 73956 6016 73958
rect 6040 73956 6096 73958
rect 36520 74010 36576 74012
rect 36600 74010 36656 74012
rect 36680 74010 36736 74012
rect 36760 74010 36816 74012
rect 36520 73958 36566 74010
rect 36566 73958 36576 74010
rect 36600 73958 36630 74010
rect 36630 73958 36642 74010
rect 36642 73958 36656 74010
rect 36680 73958 36694 74010
rect 36694 73958 36706 74010
rect 36706 73958 36736 74010
rect 36760 73958 36770 74010
rect 36770 73958 36816 74010
rect 36520 73956 36576 73958
rect 36600 73956 36656 73958
rect 36680 73956 36736 73958
rect 36760 73956 36816 73958
rect 67240 74010 67296 74012
rect 67320 74010 67376 74012
rect 67400 74010 67456 74012
rect 67480 74010 67536 74012
rect 67240 73958 67286 74010
rect 67286 73958 67296 74010
rect 67320 73958 67350 74010
rect 67350 73958 67362 74010
rect 67362 73958 67376 74010
rect 67400 73958 67414 74010
rect 67414 73958 67426 74010
rect 67426 73958 67456 74010
rect 67480 73958 67490 74010
rect 67490 73958 67536 74010
rect 67240 73956 67296 73958
rect 67320 73956 67376 73958
rect 67400 73956 67456 73958
rect 67480 73956 67536 73958
rect 5140 73466 5196 73468
rect 5220 73466 5276 73468
rect 5300 73466 5356 73468
rect 5380 73466 5436 73468
rect 5140 73414 5186 73466
rect 5186 73414 5196 73466
rect 5220 73414 5250 73466
rect 5250 73414 5262 73466
rect 5262 73414 5276 73466
rect 5300 73414 5314 73466
rect 5314 73414 5326 73466
rect 5326 73414 5356 73466
rect 5380 73414 5390 73466
rect 5390 73414 5436 73466
rect 5140 73412 5196 73414
rect 5220 73412 5276 73414
rect 5300 73412 5356 73414
rect 5380 73412 5436 73414
rect 35860 73466 35916 73468
rect 35940 73466 35996 73468
rect 36020 73466 36076 73468
rect 36100 73466 36156 73468
rect 35860 73414 35906 73466
rect 35906 73414 35916 73466
rect 35940 73414 35970 73466
rect 35970 73414 35982 73466
rect 35982 73414 35996 73466
rect 36020 73414 36034 73466
rect 36034 73414 36046 73466
rect 36046 73414 36076 73466
rect 36100 73414 36110 73466
rect 36110 73414 36156 73466
rect 35860 73412 35916 73414
rect 35940 73412 35996 73414
rect 36020 73412 36076 73414
rect 36100 73412 36156 73414
rect 66580 73466 66636 73468
rect 66660 73466 66716 73468
rect 66740 73466 66796 73468
rect 66820 73466 66876 73468
rect 66580 73414 66626 73466
rect 66626 73414 66636 73466
rect 66660 73414 66690 73466
rect 66690 73414 66702 73466
rect 66702 73414 66716 73466
rect 66740 73414 66754 73466
rect 66754 73414 66766 73466
rect 66766 73414 66796 73466
rect 66820 73414 66830 73466
rect 66830 73414 66876 73466
rect 66580 73412 66636 73414
rect 66660 73412 66716 73414
rect 66740 73412 66796 73414
rect 66820 73412 66876 73414
rect 5800 72922 5856 72924
rect 5880 72922 5936 72924
rect 5960 72922 6016 72924
rect 6040 72922 6096 72924
rect 5800 72870 5846 72922
rect 5846 72870 5856 72922
rect 5880 72870 5910 72922
rect 5910 72870 5922 72922
rect 5922 72870 5936 72922
rect 5960 72870 5974 72922
rect 5974 72870 5986 72922
rect 5986 72870 6016 72922
rect 6040 72870 6050 72922
rect 6050 72870 6096 72922
rect 5800 72868 5856 72870
rect 5880 72868 5936 72870
rect 5960 72868 6016 72870
rect 6040 72868 6096 72870
rect 36520 72922 36576 72924
rect 36600 72922 36656 72924
rect 36680 72922 36736 72924
rect 36760 72922 36816 72924
rect 36520 72870 36566 72922
rect 36566 72870 36576 72922
rect 36600 72870 36630 72922
rect 36630 72870 36642 72922
rect 36642 72870 36656 72922
rect 36680 72870 36694 72922
rect 36694 72870 36706 72922
rect 36706 72870 36736 72922
rect 36760 72870 36770 72922
rect 36770 72870 36816 72922
rect 36520 72868 36576 72870
rect 36600 72868 36656 72870
rect 36680 72868 36736 72870
rect 36760 72868 36816 72870
rect 67240 72922 67296 72924
rect 67320 72922 67376 72924
rect 67400 72922 67456 72924
rect 67480 72922 67536 72924
rect 67240 72870 67286 72922
rect 67286 72870 67296 72922
rect 67320 72870 67350 72922
rect 67350 72870 67362 72922
rect 67362 72870 67376 72922
rect 67400 72870 67414 72922
rect 67414 72870 67426 72922
rect 67426 72870 67456 72922
rect 67480 72870 67490 72922
rect 67490 72870 67536 72922
rect 67240 72868 67296 72870
rect 67320 72868 67376 72870
rect 67400 72868 67456 72870
rect 67480 72868 67536 72870
rect 5140 72378 5196 72380
rect 5220 72378 5276 72380
rect 5300 72378 5356 72380
rect 5380 72378 5436 72380
rect 5140 72326 5186 72378
rect 5186 72326 5196 72378
rect 5220 72326 5250 72378
rect 5250 72326 5262 72378
rect 5262 72326 5276 72378
rect 5300 72326 5314 72378
rect 5314 72326 5326 72378
rect 5326 72326 5356 72378
rect 5380 72326 5390 72378
rect 5390 72326 5436 72378
rect 5140 72324 5196 72326
rect 5220 72324 5276 72326
rect 5300 72324 5356 72326
rect 5380 72324 5436 72326
rect 35860 72378 35916 72380
rect 35940 72378 35996 72380
rect 36020 72378 36076 72380
rect 36100 72378 36156 72380
rect 35860 72326 35906 72378
rect 35906 72326 35916 72378
rect 35940 72326 35970 72378
rect 35970 72326 35982 72378
rect 35982 72326 35996 72378
rect 36020 72326 36034 72378
rect 36034 72326 36046 72378
rect 36046 72326 36076 72378
rect 36100 72326 36110 72378
rect 36110 72326 36156 72378
rect 35860 72324 35916 72326
rect 35940 72324 35996 72326
rect 36020 72324 36076 72326
rect 36100 72324 36156 72326
rect 66580 72378 66636 72380
rect 66660 72378 66716 72380
rect 66740 72378 66796 72380
rect 66820 72378 66876 72380
rect 66580 72326 66626 72378
rect 66626 72326 66636 72378
rect 66660 72326 66690 72378
rect 66690 72326 66702 72378
rect 66702 72326 66716 72378
rect 66740 72326 66754 72378
rect 66754 72326 66766 72378
rect 66766 72326 66796 72378
rect 66820 72326 66830 72378
rect 66830 72326 66876 72378
rect 66580 72324 66636 72326
rect 66660 72324 66716 72326
rect 66740 72324 66796 72326
rect 66820 72324 66876 72326
rect 5800 71834 5856 71836
rect 5880 71834 5936 71836
rect 5960 71834 6016 71836
rect 6040 71834 6096 71836
rect 5800 71782 5846 71834
rect 5846 71782 5856 71834
rect 5880 71782 5910 71834
rect 5910 71782 5922 71834
rect 5922 71782 5936 71834
rect 5960 71782 5974 71834
rect 5974 71782 5986 71834
rect 5986 71782 6016 71834
rect 6040 71782 6050 71834
rect 6050 71782 6096 71834
rect 5800 71780 5856 71782
rect 5880 71780 5936 71782
rect 5960 71780 6016 71782
rect 6040 71780 6096 71782
rect 36520 71834 36576 71836
rect 36600 71834 36656 71836
rect 36680 71834 36736 71836
rect 36760 71834 36816 71836
rect 36520 71782 36566 71834
rect 36566 71782 36576 71834
rect 36600 71782 36630 71834
rect 36630 71782 36642 71834
rect 36642 71782 36656 71834
rect 36680 71782 36694 71834
rect 36694 71782 36706 71834
rect 36706 71782 36736 71834
rect 36760 71782 36770 71834
rect 36770 71782 36816 71834
rect 36520 71780 36576 71782
rect 36600 71780 36656 71782
rect 36680 71780 36736 71782
rect 36760 71780 36816 71782
rect 67240 71834 67296 71836
rect 67320 71834 67376 71836
rect 67400 71834 67456 71836
rect 67480 71834 67536 71836
rect 67240 71782 67286 71834
rect 67286 71782 67296 71834
rect 67320 71782 67350 71834
rect 67350 71782 67362 71834
rect 67362 71782 67376 71834
rect 67400 71782 67414 71834
rect 67414 71782 67426 71834
rect 67426 71782 67456 71834
rect 67480 71782 67490 71834
rect 67490 71782 67536 71834
rect 67240 71780 67296 71782
rect 67320 71780 67376 71782
rect 67400 71780 67456 71782
rect 67480 71780 67536 71782
rect 5140 71290 5196 71292
rect 5220 71290 5276 71292
rect 5300 71290 5356 71292
rect 5380 71290 5436 71292
rect 5140 71238 5186 71290
rect 5186 71238 5196 71290
rect 5220 71238 5250 71290
rect 5250 71238 5262 71290
rect 5262 71238 5276 71290
rect 5300 71238 5314 71290
rect 5314 71238 5326 71290
rect 5326 71238 5356 71290
rect 5380 71238 5390 71290
rect 5390 71238 5436 71290
rect 5140 71236 5196 71238
rect 5220 71236 5276 71238
rect 5300 71236 5356 71238
rect 5380 71236 5436 71238
rect 35860 71290 35916 71292
rect 35940 71290 35996 71292
rect 36020 71290 36076 71292
rect 36100 71290 36156 71292
rect 35860 71238 35906 71290
rect 35906 71238 35916 71290
rect 35940 71238 35970 71290
rect 35970 71238 35982 71290
rect 35982 71238 35996 71290
rect 36020 71238 36034 71290
rect 36034 71238 36046 71290
rect 36046 71238 36076 71290
rect 36100 71238 36110 71290
rect 36110 71238 36156 71290
rect 35860 71236 35916 71238
rect 35940 71236 35996 71238
rect 36020 71236 36076 71238
rect 36100 71236 36156 71238
rect 66580 71290 66636 71292
rect 66660 71290 66716 71292
rect 66740 71290 66796 71292
rect 66820 71290 66876 71292
rect 66580 71238 66626 71290
rect 66626 71238 66636 71290
rect 66660 71238 66690 71290
rect 66690 71238 66702 71290
rect 66702 71238 66716 71290
rect 66740 71238 66754 71290
rect 66754 71238 66766 71290
rect 66766 71238 66796 71290
rect 66820 71238 66830 71290
rect 66830 71238 66876 71290
rect 66580 71236 66636 71238
rect 66660 71236 66716 71238
rect 66740 71236 66796 71238
rect 66820 71236 66876 71238
rect 5800 70746 5856 70748
rect 5880 70746 5936 70748
rect 5960 70746 6016 70748
rect 6040 70746 6096 70748
rect 5800 70694 5846 70746
rect 5846 70694 5856 70746
rect 5880 70694 5910 70746
rect 5910 70694 5922 70746
rect 5922 70694 5936 70746
rect 5960 70694 5974 70746
rect 5974 70694 5986 70746
rect 5986 70694 6016 70746
rect 6040 70694 6050 70746
rect 6050 70694 6096 70746
rect 5800 70692 5856 70694
rect 5880 70692 5936 70694
rect 5960 70692 6016 70694
rect 6040 70692 6096 70694
rect 36520 70746 36576 70748
rect 36600 70746 36656 70748
rect 36680 70746 36736 70748
rect 36760 70746 36816 70748
rect 36520 70694 36566 70746
rect 36566 70694 36576 70746
rect 36600 70694 36630 70746
rect 36630 70694 36642 70746
rect 36642 70694 36656 70746
rect 36680 70694 36694 70746
rect 36694 70694 36706 70746
rect 36706 70694 36736 70746
rect 36760 70694 36770 70746
rect 36770 70694 36816 70746
rect 36520 70692 36576 70694
rect 36600 70692 36656 70694
rect 36680 70692 36736 70694
rect 36760 70692 36816 70694
rect 67240 70746 67296 70748
rect 67320 70746 67376 70748
rect 67400 70746 67456 70748
rect 67480 70746 67536 70748
rect 67240 70694 67286 70746
rect 67286 70694 67296 70746
rect 67320 70694 67350 70746
rect 67350 70694 67362 70746
rect 67362 70694 67376 70746
rect 67400 70694 67414 70746
rect 67414 70694 67426 70746
rect 67426 70694 67456 70746
rect 67480 70694 67490 70746
rect 67490 70694 67536 70746
rect 67240 70692 67296 70694
rect 67320 70692 67376 70694
rect 67400 70692 67456 70694
rect 67480 70692 67536 70694
rect 5140 70202 5196 70204
rect 5220 70202 5276 70204
rect 5300 70202 5356 70204
rect 5380 70202 5436 70204
rect 5140 70150 5186 70202
rect 5186 70150 5196 70202
rect 5220 70150 5250 70202
rect 5250 70150 5262 70202
rect 5262 70150 5276 70202
rect 5300 70150 5314 70202
rect 5314 70150 5326 70202
rect 5326 70150 5356 70202
rect 5380 70150 5390 70202
rect 5390 70150 5436 70202
rect 5140 70148 5196 70150
rect 5220 70148 5276 70150
rect 5300 70148 5356 70150
rect 5380 70148 5436 70150
rect 35860 70202 35916 70204
rect 35940 70202 35996 70204
rect 36020 70202 36076 70204
rect 36100 70202 36156 70204
rect 35860 70150 35906 70202
rect 35906 70150 35916 70202
rect 35940 70150 35970 70202
rect 35970 70150 35982 70202
rect 35982 70150 35996 70202
rect 36020 70150 36034 70202
rect 36034 70150 36046 70202
rect 36046 70150 36076 70202
rect 36100 70150 36110 70202
rect 36110 70150 36156 70202
rect 35860 70148 35916 70150
rect 35940 70148 35996 70150
rect 36020 70148 36076 70150
rect 36100 70148 36156 70150
rect 66580 70202 66636 70204
rect 66660 70202 66716 70204
rect 66740 70202 66796 70204
rect 66820 70202 66876 70204
rect 66580 70150 66626 70202
rect 66626 70150 66636 70202
rect 66660 70150 66690 70202
rect 66690 70150 66702 70202
rect 66702 70150 66716 70202
rect 66740 70150 66754 70202
rect 66754 70150 66766 70202
rect 66766 70150 66796 70202
rect 66820 70150 66830 70202
rect 66830 70150 66876 70202
rect 66580 70148 66636 70150
rect 66660 70148 66716 70150
rect 66740 70148 66796 70150
rect 66820 70148 66876 70150
rect 5800 69658 5856 69660
rect 5880 69658 5936 69660
rect 5960 69658 6016 69660
rect 6040 69658 6096 69660
rect 5800 69606 5846 69658
rect 5846 69606 5856 69658
rect 5880 69606 5910 69658
rect 5910 69606 5922 69658
rect 5922 69606 5936 69658
rect 5960 69606 5974 69658
rect 5974 69606 5986 69658
rect 5986 69606 6016 69658
rect 6040 69606 6050 69658
rect 6050 69606 6096 69658
rect 5800 69604 5856 69606
rect 5880 69604 5936 69606
rect 5960 69604 6016 69606
rect 6040 69604 6096 69606
rect 36520 69658 36576 69660
rect 36600 69658 36656 69660
rect 36680 69658 36736 69660
rect 36760 69658 36816 69660
rect 36520 69606 36566 69658
rect 36566 69606 36576 69658
rect 36600 69606 36630 69658
rect 36630 69606 36642 69658
rect 36642 69606 36656 69658
rect 36680 69606 36694 69658
rect 36694 69606 36706 69658
rect 36706 69606 36736 69658
rect 36760 69606 36770 69658
rect 36770 69606 36816 69658
rect 36520 69604 36576 69606
rect 36600 69604 36656 69606
rect 36680 69604 36736 69606
rect 36760 69604 36816 69606
rect 67240 69658 67296 69660
rect 67320 69658 67376 69660
rect 67400 69658 67456 69660
rect 67480 69658 67536 69660
rect 67240 69606 67286 69658
rect 67286 69606 67296 69658
rect 67320 69606 67350 69658
rect 67350 69606 67362 69658
rect 67362 69606 67376 69658
rect 67400 69606 67414 69658
rect 67414 69606 67426 69658
rect 67426 69606 67456 69658
rect 67480 69606 67490 69658
rect 67490 69606 67536 69658
rect 67240 69604 67296 69606
rect 67320 69604 67376 69606
rect 67400 69604 67456 69606
rect 67480 69604 67536 69606
rect 5140 69114 5196 69116
rect 5220 69114 5276 69116
rect 5300 69114 5356 69116
rect 5380 69114 5436 69116
rect 5140 69062 5186 69114
rect 5186 69062 5196 69114
rect 5220 69062 5250 69114
rect 5250 69062 5262 69114
rect 5262 69062 5276 69114
rect 5300 69062 5314 69114
rect 5314 69062 5326 69114
rect 5326 69062 5356 69114
rect 5380 69062 5390 69114
rect 5390 69062 5436 69114
rect 5140 69060 5196 69062
rect 5220 69060 5276 69062
rect 5300 69060 5356 69062
rect 5380 69060 5436 69062
rect 35860 69114 35916 69116
rect 35940 69114 35996 69116
rect 36020 69114 36076 69116
rect 36100 69114 36156 69116
rect 35860 69062 35906 69114
rect 35906 69062 35916 69114
rect 35940 69062 35970 69114
rect 35970 69062 35982 69114
rect 35982 69062 35996 69114
rect 36020 69062 36034 69114
rect 36034 69062 36046 69114
rect 36046 69062 36076 69114
rect 36100 69062 36110 69114
rect 36110 69062 36156 69114
rect 35860 69060 35916 69062
rect 35940 69060 35996 69062
rect 36020 69060 36076 69062
rect 36100 69060 36156 69062
rect 66580 69114 66636 69116
rect 66660 69114 66716 69116
rect 66740 69114 66796 69116
rect 66820 69114 66876 69116
rect 66580 69062 66626 69114
rect 66626 69062 66636 69114
rect 66660 69062 66690 69114
rect 66690 69062 66702 69114
rect 66702 69062 66716 69114
rect 66740 69062 66754 69114
rect 66754 69062 66766 69114
rect 66766 69062 66796 69114
rect 66820 69062 66830 69114
rect 66830 69062 66876 69114
rect 66580 69060 66636 69062
rect 66660 69060 66716 69062
rect 66740 69060 66796 69062
rect 66820 69060 66876 69062
rect 5800 68570 5856 68572
rect 5880 68570 5936 68572
rect 5960 68570 6016 68572
rect 6040 68570 6096 68572
rect 5800 68518 5846 68570
rect 5846 68518 5856 68570
rect 5880 68518 5910 68570
rect 5910 68518 5922 68570
rect 5922 68518 5936 68570
rect 5960 68518 5974 68570
rect 5974 68518 5986 68570
rect 5986 68518 6016 68570
rect 6040 68518 6050 68570
rect 6050 68518 6096 68570
rect 5800 68516 5856 68518
rect 5880 68516 5936 68518
rect 5960 68516 6016 68518
rect 6040 68516 6096 68518
rect 36520 68570 36576 68572
rect 36600 68570 36656 68572
rect 36680 68570 36736 68572
rect 36760 68570 36816 68572
rect 36520 68518 36566 68570
rect 36566 68518 36576 68570
rect 36600 68518 36630 68570
rect 36630 68518 36642 68570
rect 36642 68518 36656 68570
rect 36680 68518 36694 68570
rect 36694 68518 36706 68570
rect 36706 68518 36736 68570
rect 36760 68518 36770 68570
rect 36770 68518 36816 68570
rect 36520 68516 36576 68518
rect 36600 68516 36656 68518
rect 36680 68516 36736 68518
rect 36760 68516 36816 68518
rect 67240 68570 67296 68572
rect 67320 68570 67376 68572
rect 67400 68570 67456 68572
rect 67480 68570 67536 68572
rect 67240 68518 67286 68570
rect 67286 68518 67296 68570
rect 67320 68518 67350 68570
rect 67350 68518 67362 68570
rect 67362 68518 67376 68570
rect 67400 68518 67414 68570
rect 67414 68518 67426 68570
rect 67426 68518 67456 68570
rect 67480 68518 67490 68570
rect 67490 68518 67536 68570
rect 67240 68516 67296 68518
rect 67320 68516 67376 68518
rect 67400 68516 67456 68518
rect 67480 68516 67536 68518
rect 5140 68026 5196 68028
rect 5220 68026 5276 68028
rect 5300 68026 5356 68028
rect 5380 68026 5436 68028
rect 5140 67974 5186 68026
rect 5186 67974 5196 68026
rect 5220 67974 5250 68026
rect 5250 67974 5262 68026
rect 5262 67974 5276 68026
rect 5300 67974 5314 68026
rect 5314 67974 5326 68026
rect 5326 67974 5356 68026
rect 5380 67974 5390 68026
rect 5390 67974 5436 68026
rect 5140 67972 5196 67974
rect 5220 67972 5276 67974
rect 5300 67972 5356 67974
rect 5380 67972 5436 67974
rect 35860 68026 35916 68028
rect 35940 68026 35996 68028
rect 36020 68026 36076 68028
rect 36100 68026 36156 68028
rect 35860 67974 35906 68026
rect 35906 67974 35916 68026
rect 35940 67974 35970 68026
rect 35970 67974 35982 68026
rect 35982 67974 35996 68026
rect 36020 67974 36034 68026
rect 36034 67974 36046 68026
rect 36046 67974 36076 68026
rect 36100 67974 36110 68026
rect 36110 67974 36156 68026
rect 35860 67972 35916 67974
rect 35940 67972 35996 67974
rect 36020 67972 36076 67974
rect 36100 67972 36156 67974
rect 66580 68026 66636 68028
rect 66660 68026 66716 68028
rect 66740 68026 66796 68028
rect 66820 68026 66876 68028
rect 66580 67974 66626 68026
rect 66626 67974 66636 68026
rect 66660 67974 66690 68026
rect 66690 67974 66702 68026
rect 66702 67974 66716 68026
rect 66740 67974 66754 68026
rect 66754 67974 66766 68026
rect 66766 67974 66796 68026
rect 66820 67974 66830 68026
rect 66830 67974 66876 68026
rect 66580 67972 66636 67974
rect 66660 67972 66716 67974
rect 66740 67972 66796 67974
rect 66820 67972 66876 67974
rect 5800 67482 5856 67484
rect 5880 67482 5936 67484
rect 5960 67482 6016 67484
rect 6040 67482 6096 67484
rect 5800 67430 5846 67482
rect 5846 67430 5856 67482
rect 5880 67430 5910 67482
rect 5910 67430 5922 67482
rect 5922 67430 5936 67482
rect 5960 67430 5974 67482
rect 5974 67430 5986 67482
rect 5986 67430 6016 67482
rect 6040 67430 6050 67482
rect 6050 67430 6096 67482
rect 5800 67428 5856 67430
rect 5880 67428 5936 67430
rect 5960 67428 6016 67430
rect 6040 67428 6096 67430
rect 36520 67482 36576 67484
rect 36600 67482 36656 67484
rect 36680 67482 36736 67484
rect 36760 67482 36816 67484
rect 36520 67430 36566 67482
rect 36566 67430 36576 67482
rect 36600 67430 36630 67482
rect 36630 67430 36642 67482
rect 36642 67430 36656 67482
rect 36680 67430 36694 67482
rect 36694 67430 36706 67482
rect 36706 67430 36736 67482
rect 36760 67430 36770 67482
rect 36770 67430 36816 67482
rect 36520 67428 36576 67430
rect 36600 67428 36656 67430
rect 36680 67428 36736 67430
rect 36760 67428 36816 67430
rect 67240 67482 67296 67484
rect 67320 67482 67376 67484
rect 67400 67482 67456 67484
rect 67480 67482 67536 67484
rect 67240 67430 67286 67482
rect 67286 67430 67296 67482
rect 67320 67430 67350 67482
rect 67350 67430 67362 67482
rect 67362 67430 67376 67482
rect 67400 67430 67414 67482
rect 67414 67430 67426 67482
rect 67426 67430 67456 67482
rect 67480 67430 67490 67482
rect 67490 67430 67536 67482
rect 67240 67428 67296 67430
rect 67320 67428 67376 67430
rect 67400 67428 67456 67430
rect 67480 67428 67536 67430
rect 5140 66938 5196 66940
rect 5220 66938 5276 66940
rect 5300 66938 5356 66940
rect 5380 66938 5436 66940
rect 5140 66886 5186 66938
rect 5186 66886 5196 66938
rect 5220 66886 5250 66938
rect 5250 66886 5262 66938
rect 5262 66886 5276 66938
rect 5300 66886 5314 66938
rect 5314 66886 5326 66938
rect 5326 66886 5356 66938
rect 5380 66886 5390 66938
rect 5390 66886 5436 66938
rect 5140 66884 5196 66886
rect 5220 66884 5276 66886
rect 5300 66884 5356 66886
rect 5380 66884 5436 66886
rect 35860 66938 35916 66940
rect 35940 66938 35996 66940
rect 36020 66938 36076 66940
rect 36100 66938 36156 66940
rect 35860 66886 35906 66938
rect 35906 66886 35916 66938
rect 35940 66886 35970 66938
rect 35970 66886 35982 66938
rect 35982 66886 35996 66938
rect 36020 66886 36034 66938
rect 36034 66886 36046 66938
rect 36046 66886 36076 66938
rect 36100 66886 36110 66938
rect 36110 66886 36156 66938
rect 35860 66884 35916 66886
rect 35940 66884 35996 66886
rect 36020 66884 36076 66886
rect 36100 66884 36156 66886
rect 66580 66938 66636 66940
rect 66660 66938 66716 66940
rect 66740 66938 66796 66940
rect 66820 66938 66876 66940
rect 66580 66886 66626 66938
rect 66626 66886 66636 66938
rect 66660 66886 66690 66938
rect 66690 66886 66702 66938
rect 66702 66886 66716 66938
rect 66740 66886 66754 66938
rect 66754 66886 66766 66938
rect 66766 66886 66796 66938
rect 66820 66886 66830 66938
rect 66830 66886 66876 66938
rect 66580 66884 66636 66886
rect 66660 66884 66716 66886
rect 66740 66884 66796 66886
rect 66820 66884 66876 66886
rect 5800 66394 5856 66396
rect 5880 66394 5936 66396
rect 5960 66394 6016 66396
rect 6040 66394 6096 66396
rect 5800 66342 5846 66394
rect 5846 66342 5856 66394
rect 5880 66342 5910 66394
rect 5910 66342 5922 66394
rect 5922 66342 5936 66394
rect 5960 66342 5974 66394
rect 5974 66342 5986 66394
rect 5986 66342 6016 66394
rect 6040 66342 6050 66394
rect 6050 66342 6096 66394
rect 5800 66340 5856 66342
rect 5880 66340 5936 66342
rect 5960 66340 6016 66342
rect 6040 66340 6096 66342
rect 36520 66394 36576 66396
rect 36600 66394 36656 66396
rect 36680 66394 36736 66396
rect 36760 66394 36816 66396
rect 36520 66342 36566 66394
rect 36566 66342 36576 66394
rect 36600 66342 36630 66394
rect 36630 66342 36642 66394
rect 36642 66342 36656 66394
rect 36680 66342 36694 66394
rect 36694 66342 36706 66394
rect 36706 66342 36736 66394
rect 36760 66342 36770 66394
rect 36770 66342 36816 66394
rect 36520 66340 36576 66342
rect 36600 66340 36656 66342
rect 36680 66340 36736 66342
rect 36760 66340 36816 66342
rect 67240 66394 67296 66396
rect 67320 66394 67376 66396
rect 67400 66394 67456 66396
rect 67480 66394 67536 66396
rect 67240 66342 67286 66394
rect 67286 66342 67296 66394
rect 67320 66342 67350 66394
rect 67350 66342 67362 66394
rect 67362 66342 67376 66394
rect 67400 66342 67414 66394
rect 67414 66342 67426 66394
rect 67426 66342 67456 66394
rect 67480 66342 67490 66394
rect 67490 66342 67536 66394
rect 67240 66340 67296 66342
rect 67320 66340 67376 66342
rect 67400 66340 67456 66342
rect 67480 66340 67536 66342
rect 5140 65850 5196 65852
rect 5220 65850 5276 65852
rect 5300 65850 5356 65852
rect 5380 65850 5436 65852
rect 5140 65798 5186 65850
rect 5186 65798 5196 65850
rect 5220 65798 5250 65850
rect 5250 65798 5262 65850
rect 5262 65798 5276 65850
rect 5300 65798 5314 65850
rect 5314 65798 5326 65850
rect 5326 65798 5356 65850
rect 5380 65798 5390 65850
rect 5390 65798 5436 65850
rect 5140 65796 5196 65798
rect 5220 65796 5276 65798
rect 5300 65796 5356 65798
rect 5380 65796 5436 65798
rect 35860 65850 35916 65852
rect 35940 65850 35996 65852
rect 36020 65850 36076 65852
rect 36100 65850 36156 65852
rect 35860 65798 35906 65850
rect 35906 65798 35916 65850
rect 35940 65798 35970 65850
rect 35970 65798 35982 65850
rect 35982 65798 35996 65850
rect 36020 65798 36034 65850
rect 36034 65798 36046 65850
rect 36046 65798 36076 65850
rect 36100 65798 36110 65850
rect 36110 65798 36156 65850
rect 35860 65796 35916 65798
rect 35940 65796 35996 65798
rect 36020 65796 36076 65798
rect 36100 65796 36156 65798
rect 66580 65850 66636 65852
rect 66660 65850 66716 65852
rect 66740 65850 66796 65852
rect 66820 65850 66876 65852
rect 66580 65798 66626 65850
rect 66626 65798 66636 65850
rect 66660 65798 66690 65850
rect 66690 65798 66702 65850
rect 66702 65798 66716 65850
rect 66740 65798 66754 65850
rect 66754 65798 66766 65850
rect 66766 65798 66796 65850
rect 66820 65798 66830 65850
rect 66830 65798 66876 65850
rect 66580 65796 66636 65798
rect 66660 65796 66716 65798
rect 66740 65796 66796 65798
rect 66820 65796 66876 65798
rect 5800 65306 5856 65308
rect 5880 65306 5936 65308
rect 5960 65306 6016 65308
rect 6040 65306 6096 65308
rect 5800 65254 5846 65306
rect 5846 65254 5856 65306
rect 5880 65254 5910 65306
rect 5910 65254 5922 65306
rect 5922 65254 5936 65306
rect 5960 65254 5974 65306
rect 5974 65254 5986 65306
rect 5986 65254 6016 65306
rect 6040 65254 6050 65306
rect 6050 65254 6096 65306
rect 5800 65252 5856 65254
rect 5880 65252 5936 65254
rect 5960 65252 6016 65254
rect 6040 65252 6096 65254
rect 36520 65306 36576 65308
rect 36600 65306 36656 65308
rect 36680 65306 36736 65308
rect 36760 65306 36816 65308
rect 36520 65254 36566 65306
rect 36566 65254 36576 65306
rect 36600 65254 36630 65306
rect 36630 65254 36642 65306
rect 36642 65254 36656 65306
rect 36680 65254 36694 65306
rect 36694 65254 36706 65306
rect 36706 65254 36736 65306
rect 36760 65254 36770 65306
rect 36770 65254 36816 65306
rect 36520 65252 36576 65254
rect 36600 65252 36656 65254
rect 36680 65252 36736 65254
rect 36760 65252 36816 65254
rect 67240 65306 67296 65308
rect 67320 65306 67376 65308
rect 67400 65306 67456 65308
rect 67480 65306 67536 65308
rect 67240 65254 67286 65306
rect 67286 65254 67296 65306
rect 67320 65254 67350 65306
rect 67350 65254 67362 65306
rect 67362 65254 67376 65306
rect 67400 65254 67414 65306
rect 67414 65254 67426 65306
rect 67426 65254 67456 65306
rect 67480 65254 67490 65306
rect 67490 65254 67536 65306
rect 67240 65252 67296 65254
rect 67320 65252 67376 65254
rect 67400 65252 67456 65254
rect 67480 65252 67536 65254
rect 5140 64762 5196 64764
rect 5220 64762 5276 64764
rect 5300 64762 5356 64764
rect 5380 64762 5436 64764
rect 5140 64710 5186 64762
rect 5186 64710 5196 64762
rect 5220 64710 5250 64762
rect 5250 64710 5262 64762
rect 5262 64710 5276 64762
rect 5300 64710 5314 64762
rect 5314 64710 5326 64762
rect 5326 64710 5356 64762
rect 5380 64710 5390 64762
rect 5390 64710 5436 64762
rect 5140 64708 5196 64710
rect 5220 64708 5276 64710
rect 5300 64708 5356 64710
rect 5380 64708 5436 64710
rect 35860 64762 35916 64764
rect 35940 64762 35996 64764
rect 36020 64762 36076 64764
rect 36100 64762 36156 64764
rect 35860 64710 35906 64762
rect 35906 64710 35916 64762
rect 35940 64710 35970 64762
rect 35970 64710 35982 64762
rect 35982 64710 35996 64762
rect 36020 64710 36034 64762
rect 36034 64710 36046 64762
rect 36046 64710 36076 64762
rect 36100 64710 36110 64762
rect 36110 64710 36156 64762
rect 35860 64708 35916 64710
rect 35940 64708 35996 64710
rect 36020 64708 36076 64710
rect 36100 64708 36156 64710
rect 66580 64762 66636 64764
rect 66660 64762 66716 64764
rect 66740 64762 66796 64764
rect 66820 64762 66876 64764
rect 66580 64710 66626 64762
rect 66626 64710 66636 64762
rect 66660 64710 66690 64762
rect 66690 64710 66702 64762
rect 66702 64710 66716 64762
rect 66740 64710 66754 64762
rect 66754 64710 66766 64762
rect 66766 64710 66796 64762
rect 66820 64710 66830 64762
rect 66830 64710 66876 64762
rect 66580 64708 66636 64710
rect 66660 64708 66716 64710
rect 66740 64708 66796 64710
rect 66820 64708 66876 64710
rect 5800 64218 5856 64220
rect 5880 64218 5936 64220
rect 5960 64218 6016 64220
rect 6040 64218 6096 64220
rect 5800 64166 5846 64218
rect 5846 64166 5856 64218
rect 5880 64166 5910 64218
rect 5910 64166 5922 64218
rect 5922 64166 5936 64218
rect 5960 64166 5974 64218
rect 5974 64166 5986 64218
rect 5986 64166 6016 64218
rect 6040 64166 6050 64218
rect 6050 64166 6096 64218
rect 5800 64164 5856 64166
rect 5880 64164 5936 64166
rect 5960 64164 6016 64166
rect 6040 64164 6096 64166
rect 36520 64218 36576 64220
rect 36600 64218 36656 64220
rect 36680 64218 36736 64220
rect 36760 64218 36816 64220
rect 36520 64166 36566 64218
rect 36566 64166 36576 64218
rect 36600 64166 36630 64218
rect 36630 64166 36642 64218
rect 36642 64166 36656 64218
rect 36680 64166 36694 64218
rect 36694 64166 36706 64218
rect 36706 64166 36736 64218
rect 36760 64166 36770 64218
rect 36770 64166 36816 64218
rect 36520 64164 36576 64166
rect 36600 64164 36656 64166
rect 36680 64164 36736 64166
rect 36760 64164 36816 64166
rect 67240 64218 67296 64220
rect 67320 64218 67376 64220
rect 67400 64218 67456 64220
rect 67480 64218 67536 64220
rect 67240 64166 67286 64218
rect 67286 64166 67296 64218
rect 67320 64166 67350 64218
rect 67350 64166 67362 64218
rect 67362 64166 67376 64218
rect 67400 64166 67414 64218
rect 67414 64166 67426 64218
rect 67426 64166 67456 64218
rect 67480 64166 67490 64218
rect 67490 64166 67536 64218
rect 67240 64164 67296 64166
rect 67320 64164 67376 64166
rect 67400 64164 67456 64166
rect 67480 64164 67536 64166
rect 5140 63674 5196 63676
rect 5220 63674 5276 63676
rect 5300 63674 5356 63676
rect 5380 63674 5436 63676
rect 5140 63622 5186 63674
rect 5186 63622 5196 63674
rect 5220 63622 5250 63674
rect 5250 63622 5262 63674
rect 5262 63622 5276 63674
rect 5300 63622 5314 63674
rect 5314 63622 5326 63674
rect 5326 63622 5356 63674
rect 5380 63622 5390 63674
rect 5390 63622 5436 63674
rect 5140 63620 5196 63622
rect 5220 63620 5276 63622
rect 5300 63620 5356 63622
rect 5380 63620 5436 63622
rect 35860 63674 35916 63676
rect 35940 63674 35996 63676
rect 36020 63674 36076 63676
rect 36100 63674 36156 63676
rect 35860 63622 35906 63674
rect 35906 63622 35916 63674
rect 35940 63622 35970 63674
rect 35970 63622 35982 63674
rect 35982 63622 35996 63674
rect 36020 63622 36034 63674
rect 36034 63622 36046 63674
rect 36046 63622 36076 63674
rect 36100 63622 36110 63674
rect 36110 63622 36156 63674
rect 35860 63620 35916 63622
rect 35940 63620 35996 63622
rect 36020 63620 36076 63622
rect 36100 63620 36156 63622
rect 66580 63674 66636 63676
rect 66660 63674 66716 63676
rect 66740 63674 66796 63676
rect 66820 63674 66876 63676
rect 66580 63622 66626 63674
rect 66626 63622 66636 63674
rect 66660 63622 66690 63674
rect 66690 63622 66702 63674
rect 66702 63622 66716 63674
rect 66740 63622 66754 63674
rect 66754 63622 66766 63674
rect 66766 63622 66796 63674
rect 66820 63622 66830 63674
rect 66830 63622 66876 63674
rect 66580 63620 66636 63622
rect 66660 63620 66716 63622
rect 66740 63620 66796 63622
rect 66820 63620 66876 63622
rect 5800 63130 5856 63132
rect 5880 63130 5936 63132
rect 5960 63130 6016 63132
rect 6040 63130 6096 63132
rect 5800 63078 5846 63130
rect 5846 63078 5856 63130
rect 5880 63078 5910 63130
rect 5910 63078 5922 63130
rect 5922 63078 5936 63130
rect 5960 63078 5974 63130
rect 5974 63078 5986 63130
rect 5986 63078 6016 63130
rect 6040 63078 6050 63130
rect 6050 63078 6096 63130
rect 5800 63076 5856 63078
rect 5880 63076 5936 63078
rect 5960 63076 6016 63078
rect 6040 63076 6096 63078
rect 36520 63130 36576 63132
rect 36600 63130 36656 63132
rect 36680 63130 36736 63132
rect 36760 63130 36816 63132
rect 36520 63078 36566 63130
rect 36566 63078 36576 63130
rect 36600 63078 36630 63130
rect 36630 63078 36642 63130
rect 36642 63078 36656 63130
rect 36680 63078 36694 63130
rect 36694 63078 36706 63130
rect 36706 63078 36736 63130
rect 36760 63078 36770 63130
rect 36770 63078 36816 63130
rect 36520 63076 36576 63078
rect 36600 63076 36656 63078
rect 36680 63076 36736 63078
rect 36760 63076 36816 63078
rect 67240 63130 67296 63132
rect 67320 63130 67376 63132
rect 67400 63130 67456 63132
rect 67480 63130 67536 63132
rect 67240 63078 67286 63130
rect 67286 63078 67296 63130
rect 67320 63078 67350 63130
rect 67350 63078 67362 63130
rect 67362 63078 67376 63130
rect 67400 63078 67414 63130
rect 67414 63078 67426 63130
rect 67426 63078 67456 63130
rect 67480 63078 67490 63130
rect 67490 63078 67536 63130
rect 67240 63076 67296 63078
rect 67320 63076 67376 63078
rect 67400 63076 67456 63078
rect 67480 63076 67536 63078
rect 5140 62586 5196 62588
rect 5220 62586 5276 62588
rect 5300 62586 5356 62588
rect 5380 62586 5436 62588
rect 5140 62534 5186 62586
rect 5186 62534 5196 62586
rect 5220 62534 5250 62586
rect 5250 62534 5262 62586
rect 5262 62534 5276 62586
rect 5300 62534 5314 62586
rect 5314 62534 5326 62586
rect 5326 62534 5356 62586
rect 5380 62534 5390 62586
rect 5390 62534 5436 62586
rect 5140 62532 5196 62534
rect 5220 62532 5276 62534
rect 5300 62532 5356 62534
rect 5380 62532 5436 62534
rect 35860 62586 35916 62588
rect 35940 62586 35996 62588
rect 36020 62586 36076 62588
rect 36100 62586 36156 62588
rect 35860 62534 35906 62586
rect 35906 62534 35916 62586
rect 35940 62534 35970 62586
rect 35970 62534 35982 62586
rect 35982 62534 35996 62586
rect 36020 62534 36034 62586
rect 36034 62534 36046 62586
rect 36046 62534 36076 62586
rect 36100 62534 36110 62586
rect 36110 62534 36156 62586
rect 35860 62532 35916 62534
rect 35940 62532 35996 62534
rect 36020 62532 36076 62534
rect 36100 62532 36156 62534
rect 66580 62586 66636 62588
rect 66660 62586 66716 62588
rect 66740 62586 66796 62588
rect 66820 62586 66876 62588
rect 66580 62534 66626 62586
rect 66626 62534 66636 62586
rect 66660 62534 66690 62586
rect 66690 62534 66702 62586
rect 66702 62534 66716 62586
rect 66740 62534 66754 62586
rect 66754 62534 66766 62586
rect 66766 62534 66796 62586
rect 66820 62534 66830 62586
rect 66830 62534 66876 62586
rect 66580 62532 66636 62534
rect 66660 62532 66716 62534
rect 66740 62532 66796 62534
rect 66820 62532 66876 62534
rect 5800 62042 5856 62044
rect 5880 62042 5936 62044
rect 5960 62042 6016 62044
rect 6040 62042 6096 62044
rect 5800 61990 5846 62042
rect 5846 61990 5856 62042
rect 5880 61990 5910 62042
rect 5910 61990 5922 62042
rect 5922 61990 5936 62042
rect 5960 61990 5974 62042
rect 5974 61990 5986 62042
rect 5986 61990 6016 62042
rect 6040 61990 6050 62042
rect 6050 61990 6096 62042
rect 5800 61988 5856 61990
rect 5880 61988 5936 61990
rect 5960 61988 6016 61990
rect 6040 61988 6096 61990
rect 36520 62042 36576 62044
rect 36600 62042 36656 62044
rect 36680 62042 36736 62044
rect 36760 62042 36816 62044
rect 36520 61990 36566 62042
rect 36566 61990 36576 62042
rect 36600 61990 36630 62042
rect 36630 61990 36642 62042
rect 36642 61990 36656 62042
rect 36680 61990 36694 62042
rect 36694 61990 36706 62042
rect 36706 61990 36736 62042
rect 36760 61990 36770 62042
rect 36770 61990 36816 62042
rect 36520 61988 36576 61990
rect 36600 61988 36656 61990
rect 36680 61988 36736 61990
rect 36760 61988 36816 61990
rect 67240 62042 67296 62044
rect 67320 62042 67376 62044
rect 67400 62042 67456 62044
rect 67480 62042 67536 62044
rect 67240 61990 67286 62042
rect 67286 61990 67296 62042
rect 67320 61990 67350 62042
rect 67350 61990 67362 62042
rect 67362 61990 67376 62042
rect 67400 61990 67414 62042
rect 67414 61990 67426 62042
rect 67426 61990 67456 62042
rect 67480 61990 67490 62042
rect 67490 61990 67536 62042
rect 67240 61988 67296 61990
rect 67320 61988 67376 61990
rect 67400 61988 67456 61990
rect 67480 61988 67536 61990
rect 5140 61498 5196 61500
rect 5220 61498 5276 61500
rect 5300 61498 5356 61500
rect 5380 61498 5436 61500
rect 5140 61446 5186 61498
rect 5186 61446 5196 61498
rect 5220 61446 5250 61498
rect 5250 61446 5262 61498
rect 5262 61446 5276 61498
rect 5300 61446 5314 61498
rect 5314 61446 5326 61498
rect 5326 61446 5356 61498
rect 5380 61446 5390 61498
rect 5390 61446 5436 61498
rect 5140 61444 5196 61446
rect 5220 61444 5276 61446
rect 5300 61444 5356 61446
rect 5380 61444 5436 61446
rect 35860 61498 35916 61500
rect 35940 61498 35996 61500
rect 36020 61498 36076 61500
rect 36100 61498 36156 61500
rect 35860 61446 35906 61498
rect 35906 61446 35916 61498
rect 35940 61446 35970 61498
rect 35970 61446 35982 61498
rect 35982 61446 35996 61498
rect 36020 61446 36034 61498
rect 36034 61446 36046 61498
rect 36046 61446 36076 61498
rect 36100 61446 36110 61498
rect 36110 61446 36156 61498
rect 35860 61444 35916 61446
rect 35940 61444 35996 61446
rect 36020 61444 36076 61446
rect 36100 61444 36156 61446
rect 66580 61498 66636 61500
rect 66660 61498 66716 61500
rect 66740 61498 66796 61500
rect 66820 61498 66876 61500
rect 66580 61446 66626 61498
rect 66626 61446 66636 61498
rect 66660 61446 66690 61498
rect 66690 61446 66702 61498
rect 66702 61446 66716 61498
rect 66740 61446 66754 61498
rect 66754 61446 66766 61498
rect 66766 61446 66796 61498
rect 66820 61446 66830 61498
rect 66830 61446 66876 61498
rect 66580 61444 66636 61446
rect 66660 61444 66716 61446
rect 66740 61444 66796 61446
rect 66820 61444 66876 61446
rect 5800 60954 5856 60956
rect 5880 60954 5936 60956
rect 5960 60954 6016 60956
rect 6040 60954 6096 60956
rect 5800 60902 5846 60954
rect 5846 60902 5856 60954
rect 5880 60902 5910 60954
rect 5910 60902 5922 60954
rect 5922 60902 5936 60954
rect 5960 60902 5974 60954
rect 5974 60902 5986 60954
rect 5986 60902 6016 60954
rect 6040 60902 6050 60954
rect 6050 60902 6096 60954
rect 5800 60900 5856 60902
rect 5880 60900 5936 60902
rect 5960 60900 6016 60902
rect 6040 60900 6096 60902
rect 36520 60954 36576 60956
rect 36600 60954 36656 60956
rect 36680 60954 36736 60956
rect 36760 60954 36816 60956
rect 36520 60902 36566 60954
rect 36566 60902 36576 60954
rect 36600 60902 36630 60954
rect 36630 60902 36642 60954
rect 36642 60902 36656 60954
rect 36680 60902 36694 60954
rect 36694 60902 36706 60954
rect 36706 60902 36736 60954
rect 36760 60902 36770 60954
rect 36770 60902 36816 60954
rect 36520 60900 36576 60902
rect 36600 60900 36656 60902
rect 36680 60900 36736 60902
rect 36760 60900 36816 60902
rect 67240 60954 67296 60956
rect 67320 60954 67376 60956
rect 67400 60954 67456 60956
rect 67480 60954 67536 60956
rect 67240 60902 67286 60954
rect 67286 60902 67296 60954
rect 67320 60902 67350 60954
rect 67350 60902 67362 60954
rect 67362 60902 67376 60954
rect 67400 60902 67414 60954
rect 67414 60902 67426 60954
rect 67426 60902 67456 60954
rect 67480 60902 67490 60954
rect 67490 60902 67536 60954
rect 67240 60900 67296 60902
rect 67320 60900 67376 60902
rect 67400 60900 67456 60902
rect 67480 60900 67536 60902
rect 5140 60410 5196 60412
rect 5220 60410 5276 60412
rect 5300 60410 5356 60412
rect 5380 60410 5436 60412
rect 5140 60358 5186 60410
rect 5186 60358 5196 60410
rect 5220 60358 5250 60410
rect 5250 60358 5262 60410
rect 5262 60358 5276 60410
rect 5300 60358 5314 60410
rect 5314 60358 5326 60410
rect 5326 60358 5356 60410
rect 5380 60358 5390 60410
rect 5390 60358 5436 60410
rect 5140 60356 5196 60358
rect 5220 60356 5276 60358
rect 5300 60356 5356 60358
rect 5380 60356 5436 60358
rect 35860 60410 35916 60412
rect 35940 60410 35996 60412
rect 36020 60410 36076 60412
rect 36100 60410 36156 60412
rect 35860 60358 35906 60410
rect 35906 60358 35916 60410
rect 35940 60358 35970 60410
rect 35970 60358 35982 60410
rect 35982 60358 35996 60410
rect 36020 60358 36034 60410
rect 36034 60358 36046 60410
rect 36046 60358 36076 60410
rect 36100 60358 36110 60410
rect 36110 60358 36156 60410
rect 35860 60356 35916 60358
rect 35940 60356 35996 60358
rect 36020 60356 36076 60358
rect 36100 60356 36156 60358
rect 66580 60410 66636 60412
rect 66660 60410 66716 60412
rect 66740 60410 66796 60412
rect 66820 60410 66876 60412
rect 66580 60358 66626 60410
rect 66626 60358 66636 60410
rect 66660 60358 66690 60410
rect 66690 60358 66702 60410
rect 66702 60358 66716 60410
rect 66740 60358 66754 60410
rect 66754 60358 66766 60410
rect 66766 60358 66796 60410
rect 66820 60358 66830 60410
rect 66830 60358 66876 60410
rect 66580 60356 66636 60358
rect 66660 60356 66716 60358
rect 66740 60356 66796 60358
rect 66820 60356 66876 60358
rect 5800 59866 5856 59868
rect 5880 59866 5936 59868
rect 5960 59866 6016 59868
rect 6040 59866 6096 59868
rect 5800 59814 5846 59866
rect 5846 59814 5856 59866
rect 5880 59814 5910 59866
rect 5910 59814 5922 59866
rect 5922 59814 5936 59866
rect 5960 59814 5974 59866
rect 5974 59814 5986 59866
rect 5986 59814 6016 59866
rect 6040 59814 6050 59866
rect 6050 59814 6096 59866
rect 5800 59812 5856 59814
rect 5880 59812 5936 59814
rect 5960 59812 6016 59814
rect 6040 59812 6096 59814
rect 36520 59866 36576 59868
rect 36600 59866 36656 59868
rect 36680 59866 36736 59868
rect 36760 59866 36816 59868
rect 36520 59814 36566 59866
rect 36566 59814 36576 59866
rect 36600 59814 36630 59866
rect 36630 59814 36642 59866
rect 36642 59814 36656 59866
rect 36680 59814 36694 59866
rect 36694 59814 36706 59866
rect 36706 59814 36736 59866
rect 36760 59814 36770 59866
rect 36770 59814 36816 59866
rect 36520 59812 36576 59814
rect 36600 59812 36656 59814
rect 36680 59812 36736 59814
rect 36760 59812 36816 59814
rect 67240 59866 67296 59868
rect 67320 59866 67376 59868
rect 67400 59866 67456 59868
rect 67480 59866 67536 59868
rect 67240 59814 67286 59866
rect 67286 59814 67296 59866
rect 67320 59814 67350 59866
rect 67350 59814 67362 59866
rect 67362 59814 67376 59866
rect 67400 59814 67414 59866
rect 67414 59814 67426 59866
rect 67426 59814 67456 59866
rect 67480 59814 67490 59866
rect 67490 59814 67536 59866
rect 67240 59812 67296 59814
rect 67320 59812 67376 59814
rect 67400 59812 67456 59814
rect 67480 59812 67536 59814
rect 5140 59322 5196 59324
rect 5220 59322 5276 59324
rect 5300 59322 5356 59324
rect 5380 59322 5436 59324
rect 5140 59270 5186 59322
rect 5186 59270 5196 59322
rect 5220 59270 5250 59322
rect 5250 59270 5262 59322
rect 5262 59270 5276 59322
rect 5300 59270 5314 59322
rect 5314 59270 5326 59322
rect 5326 59270 5356 59322
rect 5380 59270 5390 59322
rect 5390 59270 5436 59322
rect 5140 59268 5196 59270
rect 5220 59268 5276 59270
rect 5300 59268 5356 59270
rect 5380 59268 5436 59270
rect 35860 59322 35916 59324
rect 35940 59322 35996 59324
rect 36020 59322 36076 59324
rect 36100 59322 36156 59324
rect 35860 59270 35906 59322
rect 35906 59270 35916 59322
rect 35940 59270 35970 59322
rect 35970 59270 35982 59322
rect 35982 59270 35996 59322
rect 36020 59270 36034 59322
rect 36034 59270 36046 59322
rect 36046 59270 36076 59322
rect 36100 59270 36110 59322
rect 36110 59270 36156 59322
rect 35860 59268 35916 59270
rect 35940 59268 35996 59270
rect 36020 59268 36076 59270
rect 36100 59268 36156 59270
rect 66580 59322 66636 59324
rect 66660 59322 66716 59324
rect 66740 59322 66796 59324
rect 66820 59322 66876 59324
rect 66580 59270 66626 59322
rect 66626 59270 66636 59322
rect 66660 59270 66690 59322
rect 66690 59270 66702 59322
rect 66702 59270 66716 59322
rect 66740 59270 66754 59322
rect 66754 59270 66766 59322
rect 66766 59270 66796 59322
rect 66820 59270 66830 59322
rect 66830 59270 66876 59322
rect 66580 59268 66636 59270
rect 66660 59268 66716 59270
rect 66740 59268 66796 59270
rect 66820 59268 66876 59270
rect 5800 58778 5856 58780
rect 5880 58778 5936 58780
rect 5960 58778 6016 58780
rect 6040 58778 6096 58780
rect 5800 58726 5846 58778
rect 5846 58726 5856 58778
rect 5880 58726 5910 58778
rect 5910 58726 5922 58778
rect 5922 58726 5936 58778
rect 5960 58726 5974 58778
rect 5974 58726 5986 58778
rect 5986 58726 6016 58778
rect 6040 58726 6050 58778
rect 6050 58726 6096 58778
rect 5800 58724 5856 58726
rect 5880 58724 5936 58726
rect 5960 58724 6016 58726
rect 6040 58724 6096 58726
rect 36520 58778 36576 58780
rect 36600 58778 36656 58780
rect 36680 58778 36736 58780
rect 36760 58778 36816 58780
rect 36520 58726 36566 58778
rect 36566 58726 36576 58778
rect 36600 58726 36630 58778
rect 36630 58726 36642 58778
rect 36642 58726 36656 58778
rect 36680 58726 36694 58778
rect 36694 58726 36706 58778
rect 36706 58726 36736 58778
rect 36760 58726 36770 58778
rect 36770 58726 36816 58778
rect 36520 58724 36576 58726
rect 36600 58724 36656 58726
rect 36680 58724 36736 58726
rect 36760 58724 36816 58726
rect 67240 58778 67296 58780
rect 67320 58778 67376 58780
rect 67400 58778 67456 58780
rect 67480 58778 67536 58780
rect 67240 58726 67286 58778
rect 67286 58726 67296 58778
rect 67320 58726 67350 58778
rect 67350 58726 67362 58778
rect 67362 58726 67376 58778
rect 67400 58726 67414 58778
rect 67414 58726 67426 58778
rect 67426 58726 67456 58778
rect 67480 58726 67490 58778
rect 67490 58726 67536 58778
rect 67240 58724 67296 58726
rect 67320 58724 67376 58726
rect 67400 58724 67456 58726
rect 67480 58724 67536 58726
rect 5140 58234 5196 58236
rect 5220 58234 5276 58236
rect 5300 58234 5356 58236
rect 5380 58234 5436 58236
rect 5140 58182 5186 58234
rect 5186 58182 5196 58234
rect 5220 58182 5250 58234
rect 5250 58182 5262 58234
rect 5262 58182 5276 58234
rect 5300 58182 5314 58234
rect 5314 58182 5326 58234
rect 5326 58182 5356 58234
rect 5380 58182 5390 58234
rect 5390 58182 5436 58234
rect 5140 58180 5196 58182
rect 5220 58180 5276 58182
rect 5300 58180 5356 58182
rect 5380 58180 5436 58182
rect 35860 58234 35916 58236
rect 35940 58234 35996 58236
rect 36020 58234 36076 58236
rect 36100 58234 36156 58236
rect 35860 58182 35906 58234
rect 35906 58182 35916 58234
rect 35940 58182 35970 58234
rect 35970 58182 35982 58234
rect 35982 58182 35996 58234
rect 36020 58182 36034 58234
rect 36034 58182 36046 58234
rect 36046 58182 36076 58234
rect 36100 58182 36110 58234
rect 36110 58182 36156 58234
rect 35860 58180 35916 58182
rect 35940 58180 35996 58182
rect 36020 58180 36076 58182
rect 36100 58180 36156 58182
rect 66580 58234 66636 58236
rect 66660 58234 66716 58236
rect 66740 58234 66796 58236
rect 66820 58234 66876 58236
rect 66580 58182 66626 58234
rect 66626 58182 66636 58234
rect 66660 58182 66690 58234
rect 66690 58182 66702 58234
rect 66702 58182 66716 58234
rect 66740 58182 66754 58234
rect 66754 58182 66766 58234
rect 66766 58182 66796 58234
rect 66820 58182 66830 58234
rect 66830 58182 66876 58234
rect 66580 58180 66636 58182
rect 66660 58180 66716 58182
rect 66740 58180 66796 58182
rect 66820 58180 66876 58182
rect 5800 57690 5856 57692
rect 5880 57690 5936 57692
rect 5960 57690 6016 57692
rect 6040 57690 6096 57692
rect 5800 57638 5846 57690
rect 5846 57638 5856 57690
rect 5880 57638 5910 57690
rect 5910 57638 5922 57690
rect 5922 57638 5936 57690
rect 5960 57638 5974 57690
rect 5974 57638 5986 57690
rect 5986 57638 6016 57690
rect 6040 57638 6050 57690
rect 6050 57638 6096 57690
rect 5800 57636 5856 57638
rect 5880 57636 5936 57638
rect 5960 57636 6016 57638
rect 6040 57636 6096 57638
rect 36520 57690 36576 57692
rect 36600 57690 36656 57692
rect 36680 57690 36736 57692
rect 36760 57690 36816 57692
rect 36520 57638 36566 57690
rect 36566 57638 36576 57690
rect 36600 57638 36630 57690
rect 36630 57638 36642 57690
rect 36642 57638 36656 57690
rect 36680 57638 36694 57690
rect 36694 57638 36706 57690
rect 36706 57638 36736 57690
rect 36760 57638 36770 57690
rect 36770 57638 36816 57690
rect 36520 57636 36576 57638
rect 36600 57636 36656 57638
rect 36680 57636 36736 57638
rect 36760 57636 36816 57638
rect 67240 57690 67296 57692
rect 67320 57690 67376 57692
rect 67400 57690 67456 57692
rect 67480 57690 67536 57692
rect 67240 57638 67286 57690
rect 67286 57638 67296 57690
rect 67320 57638 67350 57690
rect 67350 57638 67362 57690
rect 67362 57638 67376 57690
rect 67400 57638 67414 57690
rect 67414 57638 67426 57690
rect 67426 57638 67456 57690
rect 67480 57638 67490 57690
rect 67490 57638 67536 57690
rect 67240 57636 67296 57638
rect 67320 57636 67376 57638
rect 67400 57636 67456 57638
rect 67480 57636 67536 57638
rect 5140 57146 5196 57148
rect 5220 57146 5276 57148
rect 5300 57146 5356 57148
rect 5380 57146 5436 57148
rect 5140 57094 5186 57146
rect 5186 57094 5196 57146
rect 5220 57094 5250 57146
rect 5250 57094 5262 57146
rect 5262 57094 5276 57146
rect 5300 57094 5314 57146
rect 5314 57094 5326 57146
rect 5326 57094 5356 57146
rect 5380 57094 5390 57146
rect 5390 57094 5436 57146
rect 5140 57092 5196 57094
rect 5220 57092 5276 57094
rect 5300 57092 5356 57094
rect 5380 57092 5436 57094
rect 35860 57146 35916 57148
rect 35940 57146 35996 57148
rect 36020 57146 36076 57148
rect 36100 57146 36156 57148
rect 35860 57094 35906 57146
rect 35906 57094 35916 57146
rect 35940 57094 35970 57146
rect 35970 57094 35982 57146
rect 35982 57094 35996 57146
rect 36020 57094 36034 57146
rect 36034 57094 36046 57146
rect 36046 57094 36076 57146
rect 36100 57094 36110 57146
rect 36110 57094 36156 57146
rect 35860 57092 35916 57094
rect 35940 57092 35996 57094
rect 36020 57092 36076 57094
rect 36100 57092 36156 57094
rect 66580 57146 66636 57148
rect 66660 57146 66716 57148
rect 66740 57146 66796 57148
rect 66820 57146 66876 57148
rect 66580 57094 66626 57146
rect 66626 57094 66636 57146
rect 66660 57094 66690 57146
rect 66690 57094 66702 57146
rect 66702 57094 66716 57146
rect 66740 57094 66754 57146
rect 66754 57094 66766 57146
rect 66766 57094 66796 57146
rect 66820 57094 66830 57146
rect 66830 57094 66876 57146
rect 66580 57092 66636 57094
rect 66660 57092 66716 57094
rect 66740 57092 66796 57094
rect 66820 57092 66876 57094
rect 5800 56602 5856 56604
rect 5880 56602 5936 56604
rect 5960 56602 6016 56604
rect 6040 56602 6096 56604
rect 5800 56550 5846 56602
rect 5846 56550 5856 56602
rect 5880 56550 5910 56602
rect 5910 56550 5922 56602
rect 5922 56550 5936 56602
rect 5960 56550 5974 56602
rect 5974 56550 5986 56602
rect 5986 56550 6016 56602
rect 6040 56550 6050 56602
rect 6050 56550 6096 56602
rect 5800 56548 5856 56550
rect 5880 56548 5936 56550
rect 5960 56548 6016 56550
rect 6040 56548 6096 56550
rect 36520 56602 36576 56604
rect 36600 56602 36656 56604
rect 36680 56602 36736 56604
rect 36760 56602 36816 56604
rect 36520 56550 36566 56602
rect 36566 56550 36576 56602
rect 36600 56550 36630 56602
rect 36630 56550 36642 56602
rect 36642 56550 36656 56602
rect 36680 56550 36694 56602
rect 36694 56550 36706 56602
rect 36706 56550 36736 56602
rect 36760 56550 36770 56602
rect 36770 56550 36816 56602
rect 36520 56548 36576 56550
rect 36600 56548 36656 56550
rect 36680 56548 36736 56550
rect 36760 56548 36816 56550
rect 67240 56602 67296 56604
rect 67320 56602 67376 56604
rect 67400 56602 67456 56604
rect 67480 56602 67536 56604
rect 67240 56550 67286 56602
rect 67286 56550 67296 56602
rect 67320 56550 67350 56602
rect 67350 56550 67362 56602
rect 67362 56550 67376 56602
rect 67400 56550 67414 56602
rect 67414 56550 67426 56602
rect 67426 56550 67456 56602
rect 67480 56550 67490 56602
rect 67490 56550 67536 56602
rect 67240 56548 67296 56550
rect 67320 56548 67376 56550
rect 67400 56548 67456 56550
rect 67480 56548 67536 56550
rect 5140 56058 5196 56060
rect 5220 56058 5276 56060
rect 5300 56058 5356 56060
rect 5380 56058 5436 56060
rect 5140 56006 5186 56058
rect 5186 56006 5196 56058
rect 5220 56006 5250 56058
rect 5250 56006 5262 56058
rect 5262 56006 5276 56058
rect 5300 56006 5314 56058
rect 5314 56006 5326 56058
rect 5326 56006 5356 56058
rect 5380 56006 5390 56058
rect 5390 56006 5436 56058
rect 5140 56004 5196 56006
rect 5220 56004 5276 56006
rect 5300 56004 5356 56006
rect 5380 56004 5436 56006
rect 35860 56058 35916 56060
rect 35940 56058 35996 56060
rect 36020 56058 36076 56060
rect 36100 56058 36156 56060
rect 35860 56006 35906 56058
rect 35906 56006 35916 56058
rect 35940 56006 35970 56058
rect 35970 56006 35982 56058
rect 35982 56006 35996 56058
rect 36020 56006 36034 56058
rect 36034 56006 36046 56058
rect 36046 56006 36076 56058
rect 36100 56006 36110 56058
rect 36110 56006 36156 56058
rect 35860 56004 35916 56006
rect 35940 56004 35996 56006
rect 36020 56004 36076 56006
rect 36100 56004 36156 56006
rect 66580 56058 66636 56060
rect 66660 56058 66716 56060
rect 66740 56058 66796 56060
rect 66820 56058 66876 56060
rect 66580 56006 66626 56058
rect 66626 56006 66636 56058
rect 66660 56006 66690 56058
rect 66690 56006 66702 56058
rect 66702 56006 66716 56058
rect 66740 56006 66754 56058
rect 66754 56006 66766 56058
rect 66766 56006 66796 56058
rect 66820 56006 66830 56058
rect 66830 56006 66876 56058
rect 66580 56004 66636 56006
rect 66660 56004 66716 56006
rect 66740 56004 66796 56006
rect 66820 56004 66876 56006
rect 5800 55514 5856 55516
rect 5880 55514 5936 55516
rect 5960 55514 6016 55516
rect 6040 55514 6096 55516
rect 5800 55462 5846 55514
rect 5846 55462 5856 55514
rect 5880 55462 5910 55514
rect 5910 55462 5922 55514
rect 5922 55462 5936 55514
rect 5960 55462 5974 55514
rect 5974 55462 5986 55514
rect 5986 55462 6016 55514
rect 6040 55462 6050 55514
rect 6050 55462 6096 55514
rect 5800 55460 5856 55462
rect 5880 55460 5936 55462
rect 5960 55460 6016 55462
rect 6040 55460 6096 55462
rect 36520 55514 36576 55516
rect 36600 55514 36656 55516
rect 36680 55514 36736 55516
rect 36760 55514 36816 55516
rect 36520 55462 36566 55514
rect 36566 55462 36576 55514
rect 36600 55462 36630 55514
rect 36630 55462 36642 55514
rect 36642 55462 36656 55514
rect 36680 55462 36694 55514
rect 36694 55462 36706 55514
rect 36706 55462 36736 55514
rect 36760 55462 36770 55514
rect 36770 55462 36816 55514
rect 36520 55460 36576 55462
rect 36600 55460 36656 55462
rect 36680 55460 36736 55462
rect 36760 55460 36816 55462
rect 67240 55514 67296 55516
rect 67320 55514 67376 55516
rect 67400 55514 67456 55516
rect 67480 55514 67536 55516
rect 67240 55462 67286 55514
rect 67286 55462 67296 55514
rect 67320 55462 67350 55514
rect 67350 55462 67362 55514
rect 67362 55462 67376 55514
rect 67400 55462 67414 55514
rect 67414 55462 67426 55514
rect 67426 55462 67456 55514
rect 67480 55462 67490 55514
rect 67490 55462 67536 55514
rect 67240 55460 67296 55462
rect 67320 55460 67376 55462
rect 67400 55460 67456 55462
rect 67480 55460 67536 55462
rect 5140 54970 5196 54972
rect 5220 54970 5276 54972
rect 5300 54970 5356 54972
rect 5380 54970 5436 54972
rect 5140 54918 5186 54970
rect 5186 54918 5196 54970
rect 5220 54918 5250 54970
rect 5250 54918 5262 54970
rect 5262 54918 5276 54970
rect 5300 54918 5314 54970
rect 5314 54918 5326 54970
rect 5326 54918 5356 54970
rect 5380 54918 5390 54970
rect 5390 54918 5436 54970
rect 5140 54916 5196 54918
rect 5220 54916 5276 54918
rect 5300 54916 5356 54918
rect 5380 54916 5436 54918
rect 35860 54970 35916 54972
rect 35940 54970 35996 54972
rect 36020 54970 36076 54972
rect 36100 54970 36156 54972
rect 35860 54918 35906 54970
rect 35906 54918 35916 54970
rect 35940 54918 35970 54970
rect 35970 54918 35982 54970
rect 35982 54918 35996 54970
rect 36020 54918 36034 54970
rect 36034 54918 36046 54970
rect 36046 54918 36076 54970
rect 36100 54918 36110 54970
rect 36110 54918 36156 54970
rect 35860 54916 35916 54918
rect 35940 54916 35996 54918
rect 36020 54916 36076 54918
rect 36100 54916 36156 54918
rect 66580 54970 66636 54972
rect 66660 54970 66716 54972
rect 66740 54970 66796 54972
rect 66820 54970 66876 54972
rect 66580 54918 66626 54970
rect 66626 54918 66636 54970
rect 66660 54918 66690 54970
rect 66690 54918 66702 54970
rect 66702 54918 66716 54970
rect 66740 54918 66754 54970
rect 66754 54918 66766 54970
rect 66766 54918 66796 54970
rect 66820 54918 66830 54970
rect 66830 54918 66876 54970
rect 66580 54916 66636 54918
rect 66660 54916 66716 54918
rect 66740 54916 66796 54918
rect 66820 54916 66876 54918
rect 5800 54426 5856 54428
rect 5880 54426 5936 54428
rect 5960 54426 6016 54428
rect 6040 54426 6096 54428
rect 5800 54374 5846 54426
rect 5846 54374 5856 54426
rect 5880 54374 5910 54426
rect 5910 54374 5922 54426
rect 5922 54374 5936 54426
rect 5960 54374 5974 54426
rect 5974 54374 5986 54426
rect 5986 54374 6016 54426
rect 6040 54374 6050 54426
rect 6050 54374 6096 54426
rect 5800 54372 5856 54374
rect 5880 54372 5936 54374
rect 5960 54372 6016 54374
rect 6040 54372 6096 54374
rect 36520 54426 36576 54428
rect 36600 54426 36656 54428
rect 36680 54426 36736 54428
rect 36760 54426 36816 54428
rect 36520 54374 36566 54426
rect 36566 54374 36576 54426
rect 36600 54374 36630 54426
rect 36630 54374 36642 54426
rect 36642 54374 36656 54426
rect 36680 54374 36694 54426
rect 36694 54374 36706 54426
rect 36706 54374 36736 54426
rect 36760 54374 36770 54426
rect 36770 54374 36816 54426
rect 36520 54372 36576 54374
rect 36600 54372 36656 54374
rect 36680 54372 36736 54374
rect 36760 54372 36816 54374
rect 67240 54426 67296 54428
rect 67320 54426 67376 54428
rect 67400 54426 67456 54428
rect 67480 54426 67536 54428
rect 67240 54374 67286 54426
rect 67286 54374 67296 54426
rect 67320 54374 67350 54426
rect 67350 54374 67362 54426
rect 67362 54374 67376 54426
rect 67400 54374 67414 54426
rect 67414 54374 67426 54426
rect 67426 54374 67456 54426
rect 67480 54374 67490 54426
rect 67490 54374 67536 54426
rect 67240 54372 67296 54374
rect 67320 54372 67376 54374
rect 67400 54372 67456 54374
rect 67480 54372 67536 54374
rect 5140 53882 5196 53884
rect 5220 53882 5276 53884
rect 5300 53882 5356 53884
rect 5380 53882 5436 53884
rect 5140 53830 5186 53882
rect 5186 53830 5196 53882
rect 5220 53830 5250 53882
rect 5250 53830 5262 53882
rect 5262 53830 5276 53882
rect 5300 53830 5314 53882
rect 5314 53830 5326 53882
rect 5326 53830 5356 53882
rect 5380 53830 5390 53882
rect 5390 53830 5436 53882
rect 5140 53828 5196 53830
rect 5220 53828 5276 53830
rect 5300 53828 5356 53830
rect 5380 53828 5436 53830
rect 35860 53882 35916 53884
rect 35940 53882 35996 53884
rect 36020 53882 36076 53884
rect 36100 53882 36156 53884
rect 35860 53830 35906 53882
rect 35906 53830 35916 53882
rect 35940 53830 35970 53882
rect 35970 53830 35982 53882
rect 35982 53830 35996 53882
rect 36020 53830 36034 53882
rect 36034 53830 36046 53882
rect 36046 53830 36076 53882
rect 36100 53830 36110 53882
rect 36110 53830 36156 53882
rect 35860 53828 35916 53830
rect 35940 53828 35996 53830
rect 36020 53828 36076 53830
rect 36100 53828 36156 53830
rect 66580 53882 66636 53884
rect 66660 53882 66716 53884
rect 66740 53882 66796 53884
rect 66820 53882 66876 53884
rect 66580 53830 66626 53882
rect 66626 53830 66636 53882
rect 66660 53830 66690 53882
rect 66690 53830 66702 53882
rect 66702 53830 66716 53882
rect 66740 53830 66754 53882
rect 66754 53830 66766 53882
rect 66766 53830 66796 53882
rect 66820 53830 66830 53882
rect 66830 53830 66876 53882
rect 66580 53828 66636 53830
rect 66660 53828 66716 53830
rect 66740 53828 66796 53830
rect 66820 53828 66876 53830
rect 5800 53338 5856 53340
rect 5880 53338 5936 53340
rect 5960 53338 6016 53340
rect 6040 53338 6096 53340
rect 5800 53286 5846 53338
rect 5846 53286 5856 53338
rect 5880 53286 5910 53338
rect 5910 53286 5922 53338
rect 5922 53286 5936 53338
rect 5960 53286 5974 53338
rect 5974 53286 5986 53338
rect 5986 53286 6016 53338
rect 6040 53286 6050 53338
rect 6050 53286 6096 53338
rect 5800 53284 5856 53286
rect 5880 53284 5936 53286
rect 5960 53284 6016 53286
rect 6040 53284 6096 53286
rect 36520 53338 36576 53340
rect 36600 53338 36656 53340
rect 36680 53338 36736 53340
rect 36760 53338 36816 53340
rect 36520 53286 36566 53338
rect 36566 53286 36576 53338
rect 36600 53286 36630 53338
rect 36630 53286 36642 53338
rect 36642 53286 36656 53338
rect 36680 53286 36694 53338
rect 36694 53286 36706 53338
rect 36706 53286 36736 53338
rect 36760 53286 36770 53338
rect 36770 53286 36816 53338
rect 36520 53284 36576 53286
rect 36600 53284 36656 53286
rect 36680 53284 36736 53286
rect 36760 53284 36816 53286
rect 67240 53338 67296 53340
rect 67320 53338 67376 53340
rect 67400 53338 67456 53340
rect 67480 53338 67536 53340
rect 67240 53286 67286 53338
rect 67286 53286 67296 53338
rect 67320 53286 67350 53338
rect 67350 53286 67362 53338
rect 67362 53286 67376 53338
rect 67400 53286 67414 53338
rect 67414 53286 67426 53338
rect 67426 53286 67456 53338
rect 67480 53286 67490 53338
rect 67490 53286 67536 53338
rect 67240 53284 67296 53286
rect 67320 53284 67376 53286
rect 67400 53284 67456 53286
rect 67480 53284 67536 53286
rect 5140 52794 5196 52796
rect 5220 52794 5276 52796
rect 5300 52794 5356 52796
rect 5380 52794 5436 52796
rect 5140 52742 5186 52794
rect 5186 52742 5196 52794
rect 5220 52742 5250 52794
rect 5250 52742 5262 52794
rect 5262 52742 5276 52794
rect 5300 52742 5314 52794
rect 5314 52742 5326 52794
rect 5326 52742 5356 52794
rect 5380 52742 5390 52794
rect 5390 52742 5436 52794
rect 5140 52740 5196 52742
rect 5220 52740 5276 52742
rect 5300 52740 5356 52742
rect 5380 52740 5436 52742
rect 35860 52794 35916 52796
rect 35940 52794 35996 52796
rect 36020 52794 36076 52796
rect 36100 52794 36156 52796
rect 35860 52742 35906 52794
rect 35906 52742 35916 52794
rect 35940 52742 35970 52794
rect 35970 52742 35982 52794
rect 35982 52742 35996 52794
rect 36020 52742 36034 52794
rect 36034 52742 36046 52794
rect 36046 52742 36076 52794
rect 36100 52742 36110 52794
rect 36110 52742 36156 52794
rect 35860 52740 35916 52742
rect 35940 52740 35996 52742
rect 36020 52740 36076 52742
rect 36100 52740 36156 52742
rect 66580 52794 66636 52796
rect 66660 52794 66716 52796
rect 66740 52794 66796 52796
rect 66820 52794 66876 52796
rect 66580 52742 66626 52794
rect 66626 52742 66636 52794
rect 66660 52742 66690 52794
rect 66690 52742 66702 52794
rect 66702 52742 66716 52794
rect 66740 52742 66754 52794
rect 66754 52742 66766 52794
rect 66766 52742 66796 52794
rect 66820 52742 66830 52794
rect 66830 52742 66876 52794
rect 66580 52740 66636 52742
rect 66660 52740 66716 52742
rect 66740 52740 66796 52742
rect 66820 52740 66876 52742
rect 5800 52250 5856 52252
rect 5880 52250 5936 52252
rect 5960 52250 6016 52252
rect 6040 52250 6096 52252
rect 5800 52198 5846 52250
rect 5846 52198 5856 52250
rect 5880 52198 5910 52250
rect 5910 52198 5922 52250
rect 5922 52198 5936 52250
rect 5960 52198 5974 52250
rect 5974 52198 5986 52250
rect 5986 52198 6016 52250
rect 6040 52198 6050 52250
rect 6050 52198 6096 52250
rect 5800 52196 5856 52198
rect 5880 52196 5936 52198
rect 5960 52196 6016 52198
rect 6040 52196 6096 52198
rect 36520 52250 36576 52252
rect 36600 52250 36656 52252
rect 36680 52250 36736 52252
rect 36760 52250 36816 52252
rect 36520 52198 36566 52250
rect 36566 52198 36576 52250
rect 36600 52198 36630 52250
rect 36630 52198 36642 52250
rect 36642 52198 36656 52250
rect 36680 52198 36694 52250
rect 36694 52198 36706 52250
rect 36706 52198 36736 52250
rect 36760 52198 36770 52250
rect 36770 52198 36816 52250
rect 36520 52196 36576 52198
rect 36600 52196 36656 52198
rect 36680 52196 36736 52198
rect 36760 52196 36816 52198
rect 67240 52250 67296 52252
rect 67320 52250 67376 52252
rect 67400 52250 67456 52252
rect 67480 52250 67536 52252
rect 67240 52198 67286 52250
rect 67286 52198 67296 52250
rect 67320 52198 67350 52250
rect 67350 52198 67362 52250
rect 67362 52198 67376 52250
rect 67400 52198 67414 52250
rect 67414 52198 67426 52250
rect 67426 52198 67456 52250
rect 67480 52198 67490 52250
rect 67490 52198 67536 52250
rect 67240 52196 67296 52198
rect 67320 52196 67376 52198
rect 67400 52196 67456 52198
rect 67480 52196 67536 52198
rect 77574 51756 77576 51776
rect 77576 51756 77628 51776
rect 77628 51756 77630 51776
rect 77574 51720 77630 51756
rect 5140 51706 5196 51708
rect 5220 51706 5276 51708
rect 5300 51706 5356 51708
rect 5380 51706 5436 51708
rect 5140 51654 5186 51706
rect 5186 51654 5196 51706
rect 5220 51654 5250 51706
rect 5250 51654 5262 51706
rect 5262 51654 5276 51706
rect 5300 51654 5314 51706
rect 5314 51654 5326 51706
rect 5326 51654 5356 51706
rect 5380 51654 5390 51706
rect 5390 51654 5436 51706
rect 5140 51652 5196 51654
rect 5220 51652 5276 51654
rect 5300 51652 5356 51654
rect 5380 51652 5436 51654
rect 35860 51706 35916 51708
rect 35940 51706 35996 51708
rect 36020 51706 36076 51708
rect 36100 51706 36156 51708
rect 35860 51654 35906 51706
rect 35906 51654 35916 51706
rect 35940 51654 35970 51706
rect 35970 51654 35982 51706
rect 35982 51654 35996 51706
rect 36020 51654 36034 51706
rect 36034 51654 36046 51706
rect 36046 51654 36076 51706
rect 36100 51654 36110 51706
rect 36110 51654 36156 51706
rect 35860 51652 35916 51654
rect 35940 51652 35996 51654
rect 36020 51652 36076 51654
rect 36100 51652 36156 51654
rect 66580 51706 66636 51708
rect 66660 51706 66716 51708
rect 66740 51706 66796 51708
rect 66820 51706 66876 51708
rect 66580 51654 66626 51706
rect 66626 51654 66636 51706
rect 66660 51654 66690 51706
rect 66690 51654 66702 51706
rect 66702 51654 66716 51706
rect 66740 51654 66754 51706
rect 66754 51654 66766 51706
rect 66766 51654 66796 51706
rect 66820 51654 66830 51706
rect 66830 51654 66876 51706
rect 66580 51652 66636 51654
rect 66660 51652 66716 51654
rect 66740 51652 66796 51654
rect 66820 51652 66876 51654
rect 5800 51162 5856 51164
rect 5880 51162 5936 51164
rect 5960 51162 6016 51164
rect 6040 51162 6096 51164
rect 5800 51110 5846 51162
rect 5846 51110 5856 51162
rect 5880 51110 5910 51162
rect 5910 51110 5922 51162
rect 5922 51110 5936 51162
rect 5960 51110 5974 51162
rect 5974 51110 5986 51162
rect 5986 51110 6016 51162
rect 6040 51110 6050 51162
rect 6050 51110 6096 51162
rect 5800 51108 5856 51110
rect 5880 51108 5936 51110
rect 5960 51108 6016 51110
rect 6040 51108 6096 51110
rect 36520 51162 36576 51164
rect 36600 51162 36656 51164
rect 36680 51162 36736 51164
rect 36760 51162 36816 51164
rect 36520 51110 36566 51162
rect 36566 51110 36576 51162
rect 36600 51110 36630 51162
rect 36630 51110 36642 51162
rect 36642 51110 36656 51162
rect 36680 51110 36694 51162
rect 36694 51110 36706 51162
rect 36706 51110 36736 51162
rect 36760 51110 36770 51162
rect 36770 51110 36816 51162
rect 36520 51108 36576 51110
rect 36600 51108 36656 51110
rect 36680 51108 36736 51110
rect 36760 51108 36816 51110
rect 67240 51162 67296 51164
rect 67320 51162 67376 51164
rect 67400 51162 67456 51164
rect 67480 51162 67536 51164
rect 67240 51110 67286 51162
rect 67286 51110 67296 51162
rect 67320 51110 67350 51162
rect 67350 51110 67362 51162
rect 67362 51110 67376 51162
rect 67400 51110 67414 51162
rect 67414 51110 67426 51162
rect 67426 51110 67456 51162
rect 67480 51110 67490 51162
rect 67490 51110 67536 51162
rect 67240 51108 67296 51110
rect 67320 51108 67376 51110
rect 67400 51108 67456 51110
rect 67480 51108 67536 51110
rect 5140 50618 5196 50620
rect 5220 50618 5276 50620
rect 5300 50618 5356 50620
rect 5380 50618 5436 50620
rect 5140 50566 5186 50618
rect 5186 50566 5196 50618
rect 5220 50566 5250 50618
rect 5250 50566 5262 50618
rect 5262 50566 5276 50618
rect 5300 50566 5314 50618
rect 5314 50566 5326 50618
rect 5326 50566 5356 50618
rect 5380 50566 5390 50618
rect 5390 50566 5436 50618
rect 5140 50564 5196 50566
rect 5220 50564 5276 50566
rect 5300 50564 5356 50566
rect 5380 50564 5436 50566
rect 35860 50618 35916 50620
rect 35940 50618 35996 50620
rect 36020 50618 36076 50620
rect 36100 50618 36156 50620
rect 35860 50566 35906 50618
rect 35906 50566 35916 50618
rect 35940 50566 35970 50618
rect 35970 50566 35982 50618
rect 35982 50566 35996 50618
rect 36020 50566 36034 50618
rect 36034 50566 36046 50618
rect 36046 50566 36076 50618
rect 36100 50566 36110 50618
rect 36110 50566 36156 50618
rect 35860 50564 35916 50566
rect 35940 50564 35996 50566
rect 36020 50564 36076 50566
rect 36100 50564 36156 50566
rect 66580 50618 66636 50620
rect 66660 50618 66716 50620
rect 66740 50618 66796 50620
rect 66820 50618 66876 50620
rect 66580 50566 66626 50618
rect 66626 50566 66636 50618
rect 66660 50566 66690 50618
rect 66690 50566 66702 50618
rect 66702 50566 66716 50618
rect 66740 50566 66754 50618
rect 66754 50566 66766 50618
rect 66766 50566 66796 50618
rect 66820 50566 66830 50618
rect 66830 50566 66876 50618
rect 66580 50564 66636 50566
rect 66660 50564 66716 50566
rect 66740 50564 66796 50566
rect 66820 50564 66876 50566
rect 5800 50074 5856 50076
rect 5880 50074 5936 50076
rect 5960 50074 6016 50076
rect 6040 50074 6096 50076
rect 5800 50022 5846 50074
rect 5846 50022 5856 50074
rect 5880 50022 5910 50074
rect 5910 50022 5922 50074
rect 5922 50022 5936 50074
rect 5960 50022 5974 50074
rect 5974 50022 5986 50074
rect 5986 50022 6016 50074
rect 6040 50022 6050 50074
rect 6050 50022 6096 50074
rect 5800 50020 5856 50022
rect 5880 50020 5936 50022
rect 5960 50020 6016 50022
rect 6040 50020 6096 50022
rect 36520 50074 36576 50076
rect 36600 50074 36656 50076
rect 36680 50074 36736 50076
rect 36760 50074 36816 50076
rect 36520 50022 36566 50074
rect 36566 50022 36576 50074
rect 36600 50022 36630 50074
rect 36630 50022 36642 50074
rect 36642 50022 36656 50074
rect 36680 50022 36694 50074
rect 36694 50022 36706 50074
rect 36706 50022 36736 50074
rect 36760 50022 36770 50074
rect 36770 50022 36816 50074
rect 36520 50020 36576 50022
rect 36600 50020 36656 50022
rect 36680 50020 36736 50022
rect 36760 50020 36816 50022
rect 67240 50074 67296 50076
rect 67320 50074 67376 50076
rect 67400 50074 67456 50076
rect 67480 50074 67536 50076
rect 67240 50022 67286 50074
rect 67286 50022 67296 50074
rect 67320 50022 67350 50074
rect 67350 50022 67362 50074
rect 67362 50022 67376 50074
rect 67400 50022 67414 50074
rect 67414 50022 67426 50074
rect 67426 50022 67456 50074
rect 67480 50022 67490 50074
rect 67490 50022 67536 50074
rect 67240 50020 67296 50022
rect 67320 50020 67376 50022
rect 67400 50020 67456 50022
rect 67480 50020 67536 50022
rect 77574 49716 77576 49736
rect 77576 49716 77628 49736
rect 77628 49716 77630 49736
rect 77574 49680 77630 49716
rect 5140 49530 5196 49532
rect 5220 49530 5276 49532
rect 5300 49530 5356 49532
rect 5380 49530 5436 49532
rect 5140 49478 5186 49530
rect 5186 49478 5196 49530
rect 5220 49478 5250 49530
rect 5250 49478 5262 49530
rect 5262 49478 5276 49530
rect 5300 49478 5314 49530
rect 5314 49478 5326 49530
rect 5326 49478 5356 49530
rect 5380 49478 5390 49530
rect 5390 49478 5436 49530
rect 5140 49476 5196 49478
rect 5220 49476 5276 49478
rect 5300 49476 5356 49478
rect 5380 49476 5436 49478
rect 35860 49530 35916 49532
rect 35940 49530 35996 49532
rect 36020 49530 36076 49532
rect 36100 49530 36156 49532
rect 35860 49478 35906 49530
rect 35906 49478 35916 49530
rect 35940 49478 35970 49530
rect 35970 49478 35982 49530
rect 35982 49478 35996 49530
rect 36020 49478 36034 49530
rect 36034 49478 36046 49530
rect 36046 49478 36076 49530
rect 36100 49478 36110 49530
rect 36110 49478 36156 49530
rect 35860 49476 35916 49478
rect 35940 49476 35996 49478
rect 36020 49476 36076 49478
rect 36100 49476 36156 49478
rect 66580 49530 66636 49532
rect 66660 49530 66716 49532
rect 66740 49530 66796 49532
rect 66820 49530 66876 49532
rect 66580 49478 66626 49530
rect 66626 49478 66636 49530
rect 66660 49478 66690 49530
rect 66690 49478 66702 49530
rect 66702 49478 66716 49530
rect 66740 49478 66754 49530
rect 66754 49478 66766 49530
rect 66766 49478 66796 49530
rect 66820 49478 66830 49530
rect 66830 49478 66876 49530
rect 66580 49476 66636 49478
rect 66660 49476 66716 49478
rect 66740 49476 66796 49478
rect 66820 49476 66876 49478
rect 5800 48986 5856 48988
rect 5880 48986 5936 48988
rect 5960 48986 6016 48988
rect 6040 48986 6096 48988
rect 5800 48934 5846 48986
rect 5846 48934 5856 48986
rect 5880 48934 5910 48986
rect 5910 48934 5922 48986
rect 5922 48934 5936 48986
rect 5960 48934 5974 48986
rect 5974 48934 5986 48986
rect 5986 48934 6016 48986
rect 6040 48934 6050 48986
rect 6050 48934 6096 48986
rect 5800 48932 5856 48934
rect 5880 48932 5936 48934
rect 5960 48932 6016 48934
rect 6040 48932 6096 48934
rect 36520 48986 36576 48988
rect 36600 48986 36656 48988
rect 36680 48986 36736 48988
rect 36760 48986 36816 48988
rect 36520 48934 36566 48986
rect 36566 48934 36576 48986
rect 36600 48934 36630 48986
rect 36630 48934 36642 48986
rect 36642 48934 36656 48986
rect 36680 48934 36694 48986
rect 36694 48934 36706 48986
rect 36706 48934 36736 48986
rect 36760 48934 36770 48986
rect 36770 48934 36816 48986
rect 36520 48932 36576 48934
rect 36600 48932 36656 48934
rect 36680 48932 36736 48934
rect 36760 48932 36816 48934
rect 67240 48986 67296 48988
rect 67320 48986 67376 48988
rect 67400 48986 67456 48988
rect 67480 48986 67536 48988
rect 67240 48934 67286 48986
rect 67286 48934 67296 48986
rect 67320 48934 67350 48986
rect 67350 48934 67362 48986
rect 67362 48934 67376 48986
rect 67400 48934 67414 48986
rect 67414 48934 67426 48986
rect 67426 48934 67456 48986
rect 67480 48934 67490 48986
rect 67490 48934 67536 48986
rect 67240 48932 67296 48934
rect 67320 48932 67376 48934
rect 67400 48932 67456 48934
rect 67480 48932 67536 48934
rect 5140 48442 5196 48444
rect 5220 48442 5276 48444
rect 5300 48442 5356 48444
rect 5380 48442 5436 48444
rect 5140 48390 5186 48442
rect 5186 48390 5196 48442
rect 5220 48390 5250 48442
rect 5250 48390 5262 48442
rect 5262 48390 5276 48442
rect 5300 48390 5314 48442
rect 5314 48390 5326 48442
rect 5326 48390 5356 48442
rect 5380 48390 5390 48442
rect 5390 48390 5436 48442
rect 5140 48388 5196 48390
rect 5220 48388 5276 48390
rect 5300 48388 5356 48390
rect 5380 48388 5436 48390
rect 35860 48442 35916 48444
rect 35940 48442 35996 48444
rect 36020 48442 36076 48444
rect 36100 48442 36156 48444
rect 35860 48390 35906 48442
rect 35906 48390 35916 48442
rect 35940 48390 35970 48442
rect 35970 48390 35982 48442
rect 35982 48390 35996 48442
rect 36020 48390 36034 48442
rect 36034 48390 36046 48442
rect 36046 48390 36076 48442
rect 36100 48390 36110 48442
rect 36110 48390 36156 48442
rect 35860 48388 35916 48390
rect 35940 48388 35996 48390
rect 36020 48388 36076 48390
rect 36100 48388 36156 48390
rect 66580 48442 66636 48444
rect 66660 48442 66716 48444
rect 66740 48442 66796 48444
rect 66820 48442 66876 48444
rect 66580 48390 66626 48442
rect 66626 48390 66636 48442
rect 66660 48390 66690 48442
rect 66690 48390 66702 48442
rect 66702 48390 66716 48442
rect 66740 48390 66754 48442
rect 66754 48390 66766 48442
rect 66766 48390 66796 48442
rect 66820 48390 66830 48442
rect 66830 48390 66876 48442
rect 66580 48388 66636 48390
rect 66660 48388 66716 48390
rect 66740 48388 66796 48390
rect 66820 48388 66876 48390
rect 5800 47898 5856 47900
rect 5880 47898 5936 47900
rect 5960 47898 6016 47900
rect 6040 47898 6096 47900
rect 5800 47846 5846 47898
rect 5846 47846 5856 47898
rect 5880 47846 5910 47898
rect 5910 47846 5922 47898
rect 5922 47846 5936 47898
rect 5960 47846 5974 47898
rect 5974 47846 5986 47898
rect 5986 47846 6016 47898
rect 6040 47846 6050 47898
rect 6050 47846 6096 47898
rect 5800 47844 5856 47846
rect 5880 47844 5936 47846
rect 5960 47844 6016 47846
rect 6040 47844 6096 47846
rect 36520 47898 36576 47900
rect 36600 47898 36656 47900
rect 36680 47898 36736 47900
rect 36760 47898 36816 47900
rect 36520 47846 36566 47898
rect 36566 47846 36576 47898
rect 36600 47846 36630 47898
rect 36630 47846 36642 47898
rect 36642 47846 36656 47898
rect 36680 47846 36694 47898
rect 36694 47846 36706 47898
rect 36706 47846 36736 47898
rect 36760 47846 36770 47898
rect 36770 47846 36816 47898
rect 36520 47844 36576 47846
rect 36600 47844 36656 47846
rect 36680 47844 36736 47846
rect 36760 47844 36816 47846
rect 67240 47898 67296 47900
rect 67320 47898 67376 47900
rect 67400 47898 67456 47900
rect 67480 47898 67536 47900
rect 67240 47846 67286 47898
rect 67286 47846 67296 47898
rect 67320 47846 67350 47898
rect 67350 47846 67362 47898
rect 67362 47846 67376 47898
rect 67400 47846 67414 47898
rect 67414 47846 67426 47898
rect 67426 47846 67456 47898
rect 67480 47846 67490 47898
rect 67490 47846 67536 47898
rect 67240 47844 67296 47846
rect 67320 47844 67376 47846
rect 67400 47844 67456 47846
rect 67480 47844 67536 47846
rect 5140 47354 5196 47356
rect 5220 47354 5276 47356
rect 5300 47354 5356 47356
rect 5380 47354 5436 47356
rect 5140 47302 5186 47354
rect 5186 47302 5196 47354
rect 5220 47302 5250 47354
rect 5250 47302 5262 47354
rect 5262 47302 5276 47354
rect 5300 47302 5314 47354
rect 5314 47302 5326 47354
rect 5326 47302 5356 47354
rect 5380 47302 5390 47354
rect 5390 47302 5436 47354
rect 5140 47300 5196 47302
rect 5220 47300 5276 47302
rect 5300 47300 5356 47302
rect 5380 47300 5436 47302
rect 35860 47354 35916 47356
rect 35940 47354 35996 47356
rect 36020 47354 36076 47356
rect 36100 47354 36156 47356
rect 35860 47302 35906 47354
rect 35906 47302 35916 47354
rect 35940 47302 35970 47354
rect 35970 47302 35982 47354
rect 35982 47302 35996 47354
rect 36020 47302 36034 47354
rect 36034 47302 36046 47354
rect 36046 47302 36076 47354
rect 36100 47302 36110 47354
rect 36110 47302 36156 47354
rect 35860 47300 35916 47302
rect 35940 47300 35996 47302
rect 36020 47300 36076 47302
rect 36100 47300 36156 47302
rect 66580 47354 66636 47356
rect 66660 47354 66716 47356
rect 66740 47354 66796 47356
rect 66820 47354 66876 47356
rect 66580 47302 66626 47354
rect 66626 47302 66636 47354
rect 66660 47302 66690 47354
rect 66690 47302 66702 47354
rect 66702 47302 66716 47354
rect 66740 47302 66754 47354
rect 66754 47302 66766 47354
rect 66766 47302 66796 47354
rect 66820 47302 66830 47354
rect 66830 47302 66876 47354
rect 66580 47300 66636 47302
rect 66660 47300 66716 47302
rect 66740 47300 66796 47302
rect 66820 47300 66876 47302
rect 5800 46810 5856 46812
rect 5880 46810 5936 46812
rect 5960 46810 6016 46812
rect 6040 46810 6096 46812
rect 5800 46758 5846 46810
rect 5846 46758 5856 46810
rect 5880 46758 5910 46810
rect 5910 46758 5922 46810
rect 5922 46758 5936 46810
rect 5960 46758 5974 46810
rect 5974 46758 5986 46810
rect 5986 46758 6016 46810
rect 6040 46758 6050 46810
rect 6050 46758 6096 46810
rect 5800 46756 5856 46758
rect 5880 46756 5936 46758
rect 5960 46756 6016 46758
rect 6040 46756 6096 46758
rect 36520 46810 36576 46812
rect 36600 46810 36656 46812
rect 36680 46810 36736 46812
rect 36760 46810 36816 46812
rect 36520 46758 36566 46810
rect 36566 46758 36576 46810
rect 36600 46758 36630 46810
rect 36630 46758 36642 46810
rect 36642 46758 36656 46810
rect 36680 46758 36694 46810
rect 36694 46758 36706 46810
rect 36706 46758 36736 46810
rect 36760 46758 36770 46810
rect 36770 46758 36816 46810
rect 36520 46756 36576 46758
rect 36600 46756 36656 46758
rect 36680 46756 36736 46758
rect 36760 46756 36816 46758
rect 67240 46810 67296 46812
rect 67320 46810 67376 46812
rect 67400 46810 67456 46812
rect 67480 46810 67536 46812
rect 67240 46758 67286 46810
rect 67286 46758 67296 46810
rect 67320 46758 67350 46810
rect 67350 46758 67362 46810
rect 67362 46758 67376 46810
rect 67400 46758 67414 46810
rect 67414 46758 67426 46810
rect 67426 46758 67456 46810
rect 67480 46758 67490 46810
rect 67490 46758 67536 46810
rect 67240 46756 67296 46758
rect 67320 46756 67376 46758
rect 67400 46756 67456 46758
rect 67480 46756 67536 46758
rect 5140 46266 5196 46268
rect 5220 46266 5276 46268
rect 5300 46266 5356 46268
rect 5380 46266 5436 46268
rect 5140 46214 5186 46266
rect 5186 46214 5196 46266
rect 5220 46214 5250 46266
rect 5250 46214 5262 46266
rect 5262 46214 5276 46266
rect 5300 46214 5314 46266
rect 5314 46214 5326 46266
rect 5326 46214 5356 46266
rect 5380 46214 5390 46266
rect 5390 46214 5436 46266
rect 5140 46212 5196 46214
rect 5220 46212 5276 46214
rect 5300 46212 5356 46214
rect 5380 46212 5436 46214
rect 35860 46266 35916 46268
rect 35940 46266 35996 46268
rect 36020 46266 36076 46268
rect 36100 46266 36156 46268
rect 35860 46214 35906 46266
rect 35906 46214 35916 46266
rect 35940 46214 35970 46266
rect 35970 46214 35982 46266
rect 35982 46214 35996 46266
rect 36020 46214 36034 46266
rect 36034 46214 36046 46266
rect 36046 46214 36076 46266
rect 36100 46214 36110 46266
rect 36110 46214 36156 46266
rect 35860 46212 35916 46214
rect 35940 46212 35996 46214
rect 36020 46212 36076 46214
rect 36100 46212 36156 46214
rect 66580 46266 66636 46268
rect 66660 46266 66716 46268
rect 66740 46266 66796 46268
rect 66820 46266 66876 46268
rect 66580 46214 66626 46266
rect 66626 46214 66636 46266
rect 66660 46214 66690 46266
rect 66690 46214 66702 46266
rect 66702 46214 66716 46266
rect 66740 46214 66754 46266
rect 66754 46214 66766 46266
rect 66766 46214 66796 46266
rect 66820 46214 66830 46266
rect 66830 46214 66876 46266
rect 66580 46212 66636 46214
rect 66660 46212 66716 46214
rect 66740 46212 66796 46214
rect 66820 46212 66876 46214
rect 5800 45722 5856 45724
rect 5880 45722 5936 45724
rect 5960 45722 6016 45724
rect 6040 45722 6096 45724
rect 5800 45670 5846 45722
rect 5846 45670 5856 45722
rect 5880 45670 5910 45722
rect 5910 45670 5922 45722
rect 5922 45670 5936 45722
rect 5960 45670 5974 45722
rect 5974 45670 5986 45722
rect 5986 45670 6016 45722
rect 6040 45670 6050 45722
rect 6050 45670 6096 45722
rect 5800 45668 5856 45670
rect 5880 45668 5936 45670
rect 5960 45668 6016 45670
rect 6040 45668 6096 45670
rect 36520 45722 36576 45724
rect 36600 45722 36656 45724
rect 36680 45722 36736 45724
rect 36760 45722 36816 45724
rect 36520 45670 36566 45722
rect 36566 45670 36576 45722
rect 36600 45670 36630 45722
rect 36630 45670 36642 45722
rect 36642 45670 36656 45722
rect 36680 45670 36694 45722
rect 36694 45670 36706 45722
rect 36706 45670 36736 45722
rect 36760 45670 36770 45722
rect 36770 45670 36816 45722
rect 36520 45668 36576 45670
rect 36600 45668 36656 45670
rect 36680 45668 36736 45670
rect 36760 45668 36816 45670
rect 67240 45722 67296 45724
rect 67320 45722 67376 45724
rect 67400 45722 67456 45724
rect 67480 45722 67536 45724
rect 67240 45670 67286 45722
rect 67286 45670 67296 45722
rect 67320 45670 67350 45722
rect 67350 45670 67362 45722
rect 67362 45670 67376 45722
rect 67400 45670 67414 45722
rect 67414 45670 67426 45722
rect 67426 45670 67456 45722
rect 67480 45670 67490 45722
rect 67490 45670 67536 45722
rect 67240 45668 67296 45670
rect 67320 45668 67376 45670
rect 67400 45668 67456 45670
rect 67480 45668 67536 45670
rect 1306 45600 1362 45656
rect 1214 41556 1216 41576
rect 1216 41556 1268 41576
rect 1268 41556 1270 41576
rect 1214 41520 1270 41556
rect 5140 45178 5196 45180
rect 5220 45178 5276 45180
rect 5300 45178 5356 45180
rect 5380 45178 5436 45180
rect 5140 45126 5186 45178
rect 5186 45126 5196 45178
rect 5220 45126 5250 45178
rect 5250 45126 5262 45178
rect 5262 45126 5276 45178
rect 5300 45126 5314 45178
rect 5314 45126 5326 45178
rect 5326 45126 5356 45178
rect 5380 45126 5390 45178
rect 5390 45126 5436 45178
rect 5140 45124 5196 45126
rect 5220 45124 5276 45126
rect 5300 45124 5356 45126
rect 5380 45124 5436 45126
rect 35860 45178 35916 45180
rect 35940 45178 35996 45180
rect 36020 45178 36076 45180
rect 36100 45178 36156 45180
rect 35860 45126 35906 45178
rect 35906 45126 35916 45178
rect 35940 45126 35970 45178
rect 35970 45126 35982 45178
rect 35982 45126 35996 45178
rect 36020 45126 36034 45178
rect 36034 45126 36046 45178
rect 36046 45126 36076 45178
rect 36100 45126 36110 45178
rect 36110 45126 36156 45178
rect 35860 45124 35916 45126
rect 35940 45124 35996 45126
rect 36020 45124 36076 45126
rect 36100 45124 36156 45126
rect 66580 45178 66636 45180
rect 66660 45178 66716 45180
rect 66740 45178 66796 45180
rect 66820 45178 66876 45180
rect 66580 45126 66626 45178
rect 66626 45126 66636 45178
rect 66660 45126 66690 45178
rect 66690 45126 66702 45178
rect 66702 45126 66716 45178
rect 66740 45126 66754 45178
rect 66754 45126 66766 45178
rect 66766 45126 66796 45178
rect 66820 45126 66830 45178
rect 66830 45126 66876 45178
rect 66580 45124 66636 45126
rect 66660 45124 66716 45126
rect 66740 45124 66796 45126
rect 66820 45124 66876 45126
rect 5800 44634 5856 44636
rect 5880 44634 5936 44636
rect 5960 44634 6016 44636
rect 6040 44634 6096 44636
rect 5800 44582 5846 44634
rect 5846 44582 5856 44634
rect 5880 44582 5910 44634
rect 5910 44582 5922 44634
rect 5922 44582 5936 44634
rect 5960 44582 5974 44634
rect 5974 44582 5986 44634
rect 5986 44582 6016 44634
rect 6040 44582 6050 44634
rect 6050 44582 6096 44634
rect 5800 44580 5856 44582
rect 5880 44580 5936 44582
rect 5960 44580 6016 44582
rect 6040 44580 6096 44582
rect 36520 44634 36576 44636
rect 36600 44634 36656 44636
rect 36680 44634 36736 44636
rect 36760 44634 36816 44636
rect 36520 44582 36566 44634
rect 36566 44582 36576 44634
rect 36600 44582 36630 44634
rect 36630 44582 36642 44634
rect 36642 44582 36656 44634
rect 36680 44582 36694 44634
rect 36694 44582 36706 44634
rect 36706 44582 36736 44634
rect 36760 44582 36770 44634
rect 36770 44582 36816 44634
rect 36520 44580 36576 44582
rect 36600 44580 36656 44582
rect 36680 44580 36736 44582
rect 36760 44580 36816 44582
rect 67240 44634 67296 44636
rect 67320 44634 67376 44636
rect 67400 44634 67456 44636
rect 67480 44634 67536 44636
rect 67240 44582 67286 44634
rect 67286 44582 67296 44634
rect 67320 44582 67350 44634
rect 67350 44582 67362 44634
rect 67362 44582 67376 44634
rect 67400 44582 67414 44634
rect 67414 44582 67426 44634
rect 67426 44582 67456 44634
rect 67480 44582 67490 44634
rect 67490 44582 67536 44634
rect 67240 44580 67296 44582
rect 67320 44580 67376 44582
rect 67400 44580 67456 44582
rect 67480 44580 67536 44582
rect 5140 44090 5196 44092
rect 5220 44090 5276 44092
rect 5300 44090 5356 44092
rect 5380 44090 5436 44092
rect 5140 44038 5186 44090
rect 5186 44038 5196 44090
rect 5220 44038 5250 44090
rect 5250 44038 5262 44090
rect 5262 44038 5276 44090
rect 5300 44038 5314 44090
rect 5314 44038 5326 44090
rect 5326 44038 5356 44090
rect 5380 44038 5390 44090
rect 5390 44038 5436 44090
rect 5140 44036 5196 44038
rect 5220 44036 5276 44038
rect 5300 44036 5356 44038
rect 5380 44036 5436 44038
rect 35860 44090 35916 44092
rect 35940 44090 35996 44092
rect 36020 44090 36076 44092
rect 36100 44090 36156 44092
rect 35860 44038 35906 44090
rect 35906 44038 35916 44090
rect 35940 44038 35970 44090
rect 35970 44038 35982 44090
rect 35982 44038 35996 44090
rect 36020 44038 36034 44090
rect 36034 44038 36046 44090
rect 36046 44038 36076 44090
rect 36100 44038 36110 44090
rect 36110 44038 36156 44090
rect 35860 44036 35916 44038
rect 35940 44036 35996 44038
rect 36020 44036 36076 44038
rect 36100 44036 36156 44038
rect 66580 44090 66636 44092
rect 66660 44090 66716 44092
rect 66740 44090 66796 44092
rect 66820 44090 66876 44092
rect 66580 44038 66626 44090
rect 66626 44038 66636 44090
rect 66660 44038 66690 44090
rect 66690 44038 66702 44090
rect 66702 44038 66716 44090
rect 66740 44038 66754 44090
rect 66754 44038 66766 44090
rect 66766 44038 66796 44090
rect 66820 44038 66830 44090
rect 66830 44038 66876 44090
rect 66580 44036 66636 44038
rect 66660 44036 66716 44038
rect 66740 44036 66796 44038
rect 66820 44036 66876 44038
rect 5800 43546 5856 43548
rect 5880 43546 5936 43548
rect 5960 43546 6016 43548
rect 6040 43546 6096 43548
rect 5800 43494 5846 43546
rect 5846 43494 5856 43546
rect 5880 43494 5910 43546
rect 5910 43494 5922 43546
rect 5922 43494 5936 43546
rect 5960 43494 5974 43546
rect 5974 43494 5986 43546
rect 5986 43494 6016 43546
rect 6040 43494 6050 43546
rect 6050 43494 6096 43546
rect 5800 43492 5856 43494
rect 5880 43492 5936 43494
rect 5960 43492 6016 43494
rect 6040 43492 6096 43494
rect 36520 43546 36576 43548
rect 36600 43546 36656 43548
rect 36680 43546 36736 43548
rect 36760 43546 36816 43548
rect 36520 43494 36566 43546
rect 36566 43494 36576 43546
rect 36600 43494 36630 43546
rect 36630 43494 36642 43546
rect 36642 43494 36656 43546
rect 36680 43494 36694 43546
rect 36694 43494 36706 43546
rect 36706 43494 36736 43546
rect 36760 43494 36770 43546
rect 36770 43494 36816 43546
rect 36520 43492 36576 43494
rect 36600 43492 36656 43494
rect 36680 43492 36736 43494
rect 36760 43492 36816 43494
rect 5140 43002 5196 43004
rect 5220 43002 5276 43004
rect 5300 43002 5356 43004
rect 5380 43002 5436 43004
rect 5140 42950 5186 43002
rect 5186 42950 5196 43002
rect 5220 42950 5250 43002
rect 5250 42950 5262 43002
rect 5262 42950 5276 43002
rect 5300 42950 5314 43002
rect 5314 42950 5326 43002
rect 5326 42950 5356 43002
rect 5380 42950 5390 43002
rect 5390 42950 5436 43002
rect 5140 42948 5196 42950
rect 5220 42948 5276 42950
rect 5300 42948 5356 42950
rect 5380 42948 5436 42950
rect 35860 43002 35916 43004
rect 35940 43002 35996 43004
rect 36020 43002 36076 43004
rect 36100 43002 36156 43004
rect 35860 42950 35906 43002
rect 35906 42950 35916 43002
rect 35940 42950 35970 43002
rect 35970 42950 35982 43002
rect 35982 42950 35996 43002
rect 36020 42950 36034 43002
rect 36034 42950 36046 43002
rect 36046 42950 36076 43002
rect 36100 42950 36110 43002
rect 36110 42950 36156 43002
rect 35860 42948 35916 42950
rect 35940 42948 35996 42950
rect 36020 42948 36076 42950
rect 36100 42948 36156 42950
rect 5800 42458 5856 42460
rect 5880 42458 5936 42460
rect 5960 42458 6016 42460
rect 6040 42458 6096 42460
rect 5800 42406 5846 42458
rect 5846 42406 5856 42458
rect 5880 42406 5910 42458
rect 5910 42406 5922 42458
rect 5922 42406 5936 42458
rect 5960 42406 5974 42458
rect 5974 42406 5986 42458
rect 5986 42406 6016 42458
rect 6040 42406 6050 42458
rect 6050 42406 6096 42458
rect 5800 42404 5856 42406
rect 5880 42404 5936 42406
rect 5960 42404 6016 42406
rect 6040 42404 6096 42406
rect 36520 42458 36576 42460
rect 36600 42458 36656 42460
rect 36680 42458 36736 42460
rect 36760 42458 36816 42460
rect 36520 42406 36566 42458
rect 36566 42406 36576 42458
rect 36600 42406 36630 42458
rect 36630 42406 36642 42458
rect 36642 42406 36656 42458
rect 36680 42406 36694 42458
rect 36694 42406 36706 42458
rect 36706 42406 36736 42458
rect 36760 42406 36770 42458
rect 36770 42406 36816 42458
rect 36520 42404 36576 42406
rect 36600 42404 36656 42406
rect 36680 42404 36736 42406
rect 36760 42404 36816 42406
rect 5140 41914 5196 41916
rect 5220 41914 5276 41916
rect 5300 41914 5356 41916
rect 5380 41914 5436 41916
rect 5140 41862 5186 41914
rect 5186 41862 5196 41914
rect 5220 41862 5250 41914
rect 5250 41862 5262 41914
rect 5262 41862 5276 41914
rect 5300 41862 5314 41914
rect 5314 41862 5326 41914
rect 5326 41862 5356 41914
rect 5380 41862 5390 41914
rect 5390 41862 5436 41914
rect 5140 41860 5196 41862
rect 5220 41860 5276 41862
rect 5300 41860 5356 41862
rect 5380 41860 5436 41862
rect 35860 41914 35916 41916
rect 35940 41914 35996 41916
rect 36020 41914 36076 41916
rect 36100 41914 36156 41916
rect 35860 41862 35906 41914
rect 35906 41862 35916 41914
rect 35940 41862 35970 41914
rect 35970 41862 35982 41914
rect 35982 41862 35996 41914
rect 36020 41862 36034 41914
rect 36034 41862 36046 41914
rect 36046 41862 36076 41914
rect 36100 41862 36110 41914
rect 36110 41862 36156 41914
rect 35860 41860 35916 41862
rect 35940 41860 35996 41862
rect 36020 41860 36076 41862
rect 36100 41860 36156 41862
rect 5800 41370 5856 41372
rect 5880 41370 5936 41372
rect 5960 41370 6016 41372
rect 6040 41370 6096 41372
rect 5800 41318 5846 41370
rect 5846 41318 5856 41370
rect 5880 41318 5910 41370
rect 5910 41318 5922 41370
rect 5922 41318 5936 41370
rect 5960 41318 5974 41370
rect 5974 41318 5986 41370
rect 5986 41318 6016 41370
rect 6040 41318 6050 41370
rect 6050 41318 6096 41370
rect 5800 41316 5856 41318
rect 5880 41316 5936 41318
rect 5960 41316 6016 41318
rect 6040 41316 6096 41318
rect 36520 41370 36576 41372
rect 36600 41370 36656 41372
rect 36680 41370 36736 41372
rect 36760 41370 36816 41372
rect 36520 41318 36566 41370
rect 36566 41318 36576 41370
rect 36600 41318 36630 41370
rect 36630 41318 36642 41370
rect 36642 41318 36656 41370
rect 36680 41318 36694 41370
rect 36694 41318 36706 41370
rect 36706 41318 36736 41370
rect 36760 41318 36770 41370
rect 36770 41318 36816 41370
rect 36520 41316 36576 41318
rect 36600 41316 36656 41318
rect 36680 41316 36736 41318
rect 36760 41316 36816 41318
rect 5140 40826 5196 40828
rect 5220 40826 5276 40828
rect 5300 40826 5356 40828
rect 5380 40826 5436 40828
rect 5140 40774 5186 40826
rect 5186 40774 5196 40826
rect 5220 40774 5250 40826
rect 5250 40774 5262 40826
rect 5262 40774 5276 40826
rect 5300 40774 5314 40826
rect 5314 40774 5326 40826
rect 5326 40774 5356 40826
rect 5380 40774 5390 40826
rect 5390 40774 5436 40826
rect 5140 40772 5196 40774
rect 5220 40772 5276 40774
rect 5300 40772 5356 40774
rect 5380 40772 5436 40774
rect 35860 40826 35916 40828
rect 35940 40826 35996 40828
rect 36020 40826 36076 40828
rect 36100 40826 36156 40828
rect 35860 40774 35906 40826
rect 35906 40774 35916 40826
rect 35940 40774 35970 40826
rect 35970 40774 35982 40826
rect 35982 40774 35996 40826
rect 36020 40774 36034 40826
rect 36034 40774 36046 40826
rect 36046 40774 36076 40826
rect 36100 40774 36110 40826
rect 36110 40774 36156 40826
rect 35860 40772 35916 40774
rect 35940 40772 35996 40774
rect 36020 40772 36076 40774
rect 36100 40772 36156 40774
rect 5800 40282 5856 40284
rect 5880 40282 5936 40284
rect 5960 40282 6016 40284
rect 6040 40282 6096 40284
rect 5800 40230 5846 40282
rect 5846 40230 5856 40282
rect 5880 40230 5910 40282
rect 5910 40230 5922 40282
rect 5922 40230 5936 40282
rect 5960 40230 5974 40282
rect 5974 40230 5986 40282
rect 5986 40230 6016 40282
rect 6040 40230 6050 40282
rect 6050 40230 6096 40282
rect 5800 40228 5856 40230
rect 5880 40228 5936 40230
rect 5960 40228 6016 40230
rect 6040 40228 6096 40230
rect 36520 40282 36576 40284
rect 36600 40282 36656 40284
rect 36680 40282 36736 40284
rect 36760 40282 36816 40284
rect 36520 40230 36566 40282
rect 36566 40230 36576 40282
rect 36600 40230 36630 40282
rect 36630 40230 36642 40282
rect 36642 40230 36656 40282
rect 36680 40230 36694 40282
rect 36694 40230 36706 40282
rect 36706 40230 36736 40282
rect 36760 40230 36770 40282
rect 36770 40230 36816 40282
rect 36520 40228 36576 40230
rect 36600 40228 36656 40230
rect 36680 40228 36736 40230
rect 36760 40228 36816 40230
rect 5140 39738 5196 39740
rect 5220 39738 5276 39740
rect 5300 39738 5356 39740
rect 5380 39738 5436 39740
rect 5140 39686 5186 39738
rect 5186 39686 5196 39738
rect 5220 39686 5250 39738
rect 5250 39686 5262 39738
rect 5262 39686 5276 39738
rect 5300 39686 5314 39738
rect 5314 39686 5326 39738
rect 5326 39686 5356 39738
rect 5380 39686 5390 39738
rect 5390 39686 5436 39738
rect 5140 39684 5196 39686
rect 5220 39684 5276 39686
rect 5300 39684 5356 39686
rect 5380 39684 5436 39686
rect 35860 39738 35916 39740
rect 35940 39738 35996 39740
rect 36020 39738 36076 39740
rect 36100 39738 36156 39740
rect 35860 39686 35906 39738
rect 35906 39686 35916 39738
rect 35940 39686 35970 39738
rect 35970 39686 35982 39738
rect 35982 39686 35996 39738
rect 36020 39686 36034 39738
rect 36034 39686 36046 39738
rect 36046 39686 36076 39738
rect 36100 39686 36110 39738
rect 36110 39686 36156 39738
rect 35860 39684 35916 39686
rect 35940 39684 35996 39686
rect 36020 39684 36076 39686
rect 36100 39684 36156 39686
rect 5800 39194 5856 39196
rect 5880 39194 5936 39196
rect 5960 39194 6016 39196
rect 6040 39194 6096 39196
rect 5800 39142 5846 39194
rect 5846 39142 5856 39194
rect 5880 39142 5910 39194
rect 5910 39142 5922 39194
rect 5922 39142 5936 39194
rect 5960 39142 5974 39194
rect 5974 39142 5986 39194
rect 5986 39142 6016 39194
rect 6040 39142 6050 39194
rect 6050 39142 6096 39194
rect 5800 39140 5856 39142
rect 5880 39140 5936 39142
rect 5960 39140 6016 39142
rect 6040 39140 6096 39142
rect 36520 39194 36576 39196
rect 36600 39194 36656 39196
rect 36680 39194 36736 39196
rect 36760 39194 36816 39196
rect 36520 39142 36566 39194
rect 36566 39142 36576 39194
rect 36600 39142 36630 39194
rect 36630 39142 36642 39194
rect 36642 39142 36656 39194
rect 36680 39142 36694 39194
rect 36694 39142 36706 39194
rect 36706 39142 36736 39194
rect 36760 39142 36770 39194
rect 36770 39142 36816 39194
rect 36520 39140 36576 39142
rect 36600 39140 36656 39142
rect 36680 39140 36736 39142
rect 36760 39140 36816 39142
rect 5140 38650 5196 38652
rect 5220 38650 5276 38652
rect 5300 38650 5356 38652
rect 5380 38650 5436 38652
rect 5140 38598 5186 38650
rect 5186 38598 5196 38650
rect 5220 38598 5250 38650
rect 5250 38598 5262 38650
rect 5262 38598 5276 38650
rect 5300 38598 5314 38650
rect 5314 38598 5326 38650
rect 5326 38598 5356 38650
rect 5380 38598 5390 38650
rect 5390 38598 5436 38650
rect 5140 38596 5196 38598
rect 5220 38596 5276 38598
rect 5300 38596 5356 38598
rect 5380 38596 5436 38598
rect 35860 38650 35916 38652
rect 35940 38650 35996 38652
rect 36020 38650 36076 38652
rect 36100 38650 36156 38652
rect 35860 38598 35906 38650
rect 35906 38598 35916 38650
rect 35940 38598 35970 38650
rect 35970 38598 35982 38650
rect 35982 38598 35996 38650
rect 36020 38598 36034 38650
rect 36034 38598 36046 38650
rect 36046 38598 36076 38650
rect 36100 38598 36110 38650
rect 36110 38598 36156 38650
rect 35860 38596 35916 38598
rect 35940 38596 35996 38598
rect 36020 38596 36076 38598
rect 36100 38596 36156 38598
rect 5800 38106 5856 38108
rect 5880 38106 5936 38108
rect 5960 38106 6016 38108
rect 6040 38106 6096 38108
rect 5800 38054 5846 38106
rect 5846 38054 5856 38106
rect 5880 38054 5910 38106
rect 5910 38054 5922 38106
rect 5922 38054 5936 38106
rect 5960 38054 5974 38106
rect 5974 38054 5986 38106
rect 5986 38054 6016 38106
rect 6040 38054 6050 38106
rect 6050 38054 6096 38106
rect 5800 38052 5856 38054
rect 5880 38052 5936 38054
rect 5960 38052 6016 38054
rect 6040 38052 6096 38054
rect 36520 38106 36576 38108
rect 36600 38106 36656 38108
rect 36680 38106 36736 38108
rect 36760 38106 36816 38108
rect 36520 38054 36566 38106
rect 36566 38054 36576 38106
rect 36600 38054 36630 38106
rect 36630 38054 36642 38106
rect 36642 38054 36656 38106
rect 36680 38054 36694 38106
rect 36694 38054 36706 38106
rect 36706 38054 36736 38106
rect 36760 38054 36770 38106
rect 36770 38054 36816 38106
rect 36520 38052 36576 38054
rect 36600 38052 36656 38054
rect 36680 38052 36736 38054
rect 36760 38052 36816 38054
rect 5140 37562 5196 37564
rect 5220 37562 5276 37564
rect 5300 37562 5356 37564
rect 5380 37562 5436 37564
rect 5140 37510 5186 37562
rect 5186 37510 5196 37562
rect 5220 37510 5250 37562
rect 5250 37510 5262 37562
rect 5262 37510 5276 37562
rect 5300 37510 5314 37562
rect 5314 37510 5326 37562
rect 5326 37510 5356 37562
rect 5380 37510 5390 37562
rect 5390 37510 5436 37562
rect 5140 37508 5196 37510
rect 5220 37508 5276 37510
rect 5300 37508 5356 37510
rect 5380 37508 5436 37510
rect 35860 37562 35916 37564
rect 35940 37562 35996 37564
rect 36020 37562 36076 37564
rect 36100 37562 36156 37564
rect 35860 37510 35906 37562
rect 35906 37510 35916 37562
rect 35940 37510 35970 37562
rect 35970 37510 35982 37562
rect 35982 37510 35996 37562
rect 36020 37510 36034 37562
rect 36034 37510 36046 37562
rect 36046 37510 36076 37562
rect 36100 37510 36110 37562
rect 36110 37510 36156 37562
rect 35860 37508 35916 37510
rect 35940 37508 35996 37510
rect 36020 37508 36076 37510
rect 36100 37508 36156 37510
rect 5800 37018 5856 37020
rect 5880 37018 5936 37020
rect 5960 37018 6016 37020
rect 6040 37018 6096 37020
rect 5800 36966 5846 37018
rect 5846 36966 5856 37018
rect 5880 36966 5910 37018
rect 5910 36966 5922 37018
rect 5922 36966 5936 37018
rect 5960 36966 5974 37018
rect 5974 36966 5986 37018
rect 5986 36966 6016 37018
rect 6040 36966 6050 37018
rect 6050 36966 6096 37018
rect 5800 36964 5856 36966
rect 5880 36964 5936 36966
rect 5960 36964 6016 36966
rect 6040 36964 6096 36966
rect 36520 37018 36576 37020
rect 36600 37018 36656 37020
rect 36680 37018 36736 37020
rect 36760 37018 36816 37020
rect 36520 36966 36566 37018
rect 36566 36966 36576 37018
rect 36600 36966 36630 37018
rect 36630 36966 36642 37018
rect 36642 36966 36656 37018
rect 36680 36966 36694 37018
rect 36694 36966 36706 37018
rect 36706 36966 36736 37018
rect 36760 36966 36770 37018
rect 36770 36966 36816 37018
rect 36520 36964 36576 36966
rect 36600 36964 36656 36966
rect 36680 36964 36736 36966
rect 36760 36964 36816 36966
rect 5140 36474 5196 36476
rect 5220 36474 5276 36476
rect 5300 36474 5356 36476
rect 5380 36474 5436 36476
rect 5140 36422 5186 36474
rect 5186 36422 5196 36474
rect 5220 36422 5250 36474
rect 5250 36422 5262 36474
rect 5262 36422 5276 36474
rect 5300 36422 5314 36474
rect 5314 36422 5326 36474
rect 5326 36422 5356 36474
rect 5380 36422 5390 36474
rect 5390 36422 5436 36474
rect 5140 36420 5196 36422
rect 5220 36420 5276 36422
rect 5300 36420 5356 36422
rect 5380 36420 5436 36422
rect 35860 36474 35916 36476
rect 35940 36474 35996 36476
rect 36020 36474 36076 36476
rect 36100 36474 36156 36476
rect 35860 36422 35906 36474
rect 35906 36422 35916 36474
rect 35940 36422 35970 36474
rect 35970 36422 35982 36474
rect 35982 36422 35996 36474
rect 36020 36422 36034 36474
rect 36034 36422 36046 36474
rect 36046 36422 36076 36474
rect 36100 36422 36110 36474
rect 36110 36422 36156 36474
rect 35860 36420 35916 36422
rect 35940 36420 35996 36422
rect 36020 36420 36076 36422
rect 36100 36420 36156 36422
rect 5800 35930 5856 35932
rect 5880 35930 5936 35932
rect 5960 35930 6016 35932
rect 6040 35930 6096 35932
rect 5800 35878 5846 35930
rect 5846 35878 5856 35930
rect 5880 35878 5910 35930
rect 5910 35878 5922 35930
rect 5922 35878 5936 35930
rect 5960 35878 5974 35930
rect 5974 35878 5986 35930
rect 5986 35878 6016 35930
rect 6040 35878 6050 35930
rect 6050 35878 6096 35930
rect 5800 35876 5856 35878
rect 5880 35876 5936 35878
rect 5960 35876 6016 35878
rect 6040 35876 6096 35878
rect 36520 35930 36576 35932
rect 36600 35930 36656 35932
rect 36680 35930 36736 35932
rect 36760 35930 36816 35932
rect 36520 35878 36566 35930
rect 36566 35878 36576 35930
rect 36600 35878 36630 35930
rect 36630 35878 36642 35930
rect 36642 35878 36656 35930
rect 36680 35878 36694 35930
rect 36694 35878 36706 35930
rect 36706 35878 36736 35930
rect 36760 35878 36770 35930
rect 36770 35878 36816 35930
rect 36520 35876 36576 35878
rect 36600 35876 36656 35878
rect 36680 35876 36736 35878
rect 36760 35876 36816 35878
rect 1214 35436 1216 35456
rect 1216 35436 1268 35456
rect 1268 35436 1270 35456
rect 1214 35400 1270 35436
rect 5140 35386 5196 35388
rect 5220 35386 5276 35388
rect 5300 35386 5356 35388
rect 5380 35386 5436 35388
rect 5140 35334 5186 35386
rect 5186 35334 5196 35386
rect 5220 35334 5250 35386
rect 5250 35334 5262 35386
rect 5262 35334 5276 35386
rect 5300 35334 5314 35386
rect 5314 35334 5326 35386
rect 5326 35334 5356 35386
rect 5380 35334 5390 35386
rect 5390 35334 5436 35386
rect 5140 35332 5196 35334
rect 5220 35332 5276 35334
rect 5300 35332 5356 35334
rect 5380 35332 5436 35334
rect 35860 35386 35916 35388
rect 35940 35386 35996 35388
rect 36020 35386 36076 35388
rect 36100 35386 36156 35388
rect 35860 35334 35906 35386
rect 35906 35334 35916 35386
rect 35940 35334 35970 35386
rect 35970 35334 35982 35386
rect 35982 35334 35996 35386
rect 36020 35334 36034 35386
rect 36034 35334 36046 35386
rect 36046 35334 36076 35386
rect 36100 35334 36110 35386
rect 36110 35334 36156 35386
rect 35860 35332 35916 35334
rect 35940 35332 35996 35334
rect 36020 35332 36076 35334
rect 36100 35332 36156 35334
rect 67240 43546 67296 43548
rect 67320 43546 67376 43548
rect 67400 43546 67456 43548
rect 67480 43546 67536 43548
rect 67240 43494 67286 43546
rect 67286 43494 67296 43546
rect 67320 43494 67350 43546
rect 67350 43494 67362 43546
rect 67362 43494 67376 43546
rect 67400 43494 67414 43546
rect 67414 43494 67426 43546
rect 67426 43494 67456 43546
rect 67480 43494 67490 43546
rect 67490 43494 67536 43546
rect 67240 43492 67296 43494
rect 67320 43492 67376 43494
rect 67400 43492 67456 43494
rect 67480 43492 67536 43494
rect 66580 43002 66636 43004
rect 66660 43002 66716 43004
rect 66740 43002 66796 43004
rect 66820 43002 66876 43004
rect 66580 42950 66626 43002
rect 66626 42950 66636 43002
rect 66660 42950 66690 43002
rect 66690 42950 66702 43002
rect 66702 42950 66716 43002
rect 66740 42950 66754 43002
rect 66754 42950 66766 43002
rect 66766 42950 66796 43002
rect 66820 42950 66830 43002
rect 66830 42950 66876 43002
rect 66580 42948 66636 42950
rect 66660 42948 66716 42950
rect 66740 42948 66796 42950
rect 66820 42948 66876 42950
rect 66580 41914 66636 41916
rect 66660 41914 66716 41916
rect 66740 41914 66796 41916
rect 66820 41914 66876 41916
rect 66580 41862 66626 41914
rect 66626 41862 66636 41914
rect 66660 41862 66690 41914
rect 66690 41862 66702 41914
rect 66702 41862 66716 41914
rect 66740 41862 66754 41914
rect 66754 41862 66766 41914
rect 66766 41862 66796 41914
rect 66820 41862 66830 41914
rect 66830 41862 66876 41914
rect 66580 41860 66636 41862
rect 66660 41860 66716 41862
rect 66740 41860 66796 41862
rect 66820 41860 66876 41862
rect 66580 40826 66636 40828
rect 66660 40826 66716 40828
rect 66740 40826 66796 40828
rect 66820 40826 66876 40828
rect 66580 40774 66626 40826
rect 66626 40774 66636 40826
rect 66660 40774 66690 40826
rect 66690 40774 66702 40826
rect 66702 40774 66716 40826
rect 66740 40774 66754 40826
rect 66754 40774 66766 40826
rect 66766 40774 66796 40826
rect 66820 40774 66830 40826
rect 66830 40774 66876 40826
rect 66580 40772 66636 40774
rect 66660 40772 66716 40774
rect 66740 40772 66796 40774
rect 66820 40772 66876 40774
rect 66580 39738 66636 39740
rect 66660 39738 66716 39740
rect 66740 39738 66796 39740
rect 66820 39738 66876 39740
rect 66580 39686 66626 39738
rect 66626 39686 66636 39738
rect 66660 39686 66690 39738
rect 66690 39686 66702 39738
rect 66702 39686 66716 39738
rect 66740 39686 66754 39738
rect 66754 39686 66766 39738
rect 66766 39686 66796 39738
rect 66820 39686 66830 39738
rect 66830 39686 66876 39738
rect 66580 39684 66636 39686
rect 66660 39684 66716 39686
rect 66740 39684 66796 39686
rect 66820 39684 66876 39686
rect 67240 42458 67296 42460
rect 67320 42458 67376 42460
rect 67400 42458 67456 42460
rect 67480 42458 67536 42460
rect 67240 42406 67286 42458
rect 67286 42406 67296 42458
rect 67320 42406 67350 42458
rect 67350 42406 67362 42458
rect 67362 42406 67376 42458
rect 67400 42406 67414 42458
rect 67414 42406 67426 42458
rect 67426 42406 67456 42458
rect 67480 42406 67490 42458
rect 67490 42406 67536 42458
rect 67240 42404 67296 42406
rect 67320 42404 67376 42406
rect 67400 42404 67456 42406
rect 67480 42404 67536 42406
rect 67240 41370 67296 41372
rect 67320 41370 67376 41372
rect 67400 41370 67456 41372
rect 67480 41370 67536 41372
rect 67240 41318 67286 41370
rect 67286 41318 67296 41370
rect 67320 41318 67350 41370
rect 67350 41318 67362 41370
rect 67362 41318 67376 41370
rect 67400 41318 67414 41370
rect 67414 41318 67426 41370
rect 67426 41318 67456 41370
rect 67480 41318 67490 41370
rect 67490 41318 67536 41370
rect 67240 41316 67296 41318
rect 67320 41316 67376 41318
rect 67400 41316 67456 41318
rect 67480 41316 67536 41318
rect 67240 40282 67296 40284
rect 67320 40282 67376 40284
rect 67400 40282 67456 40284
rect 67480 40282 67536 40284
rect 67240 40230 67286 40282
rect 67286 40230 67296 40282
rect 67320 40230 67350 40282
rect 67350 40230 67362 40282
rect 67362 40230 67376 40282
rect 67400 40230 67414 40282
rect 67414 40230 67426 40282
rect 67426 40230 67456 40282
rect 67480 40230 67490 40282
rect 67490 40230 67536 40282
rect 67240 40228 67296 40230
rect 67320 40228 67376 40230
rect 67400 40228 67456 40230
rect 67480 40228 67536 40230
rect 66580 38650 66636 38652
rect 66660 38650 66716 38652
rect 66740 38650 66796 38652
rect 66820 38650 66876 38652
rect 66580 38598 66626 38650
rect 66626 38598 66636 38650
rect 66660 38598 66690 38650
rect 66690 38598 66702 38650
rect 66702 38598 66716 38650
rect 66740 38598 66754 38650
rect 66754 38598 66766 38650
rect 66766 38598 66796 38650
rect 66820 38598 66830 38650
rect 66830 38598 66876 38650
rect 66580 38596 66636 38598
rect 66660 38596 66716 38598
rect 66740 38596 66796 38598
rect 66820 38596 66876 38598
rect 66580 37562 66636 37564
rect 66660 37562 66716 37564
rect 66740 37562 66796 37564
rect 66820 37562 66876 37564
rect 66580 37510 66626 37562
rect 66626 37510 66636 37562
rect 66660 37510 66690 37562
rect 66690 37510 66702 37562
rect 66702 37510 66716 37562
rect 66740 37510 66754 37562
rect 66754 37510 66766 37562
rect 66766 37510 66796 37562
rect 66820 37510 66830 37562
rect 66830 37510 66876 37562
rect 66580 37508 66636 37510
rect 66660 37508 66716 37510
rect 66740 37508 66796 37510
rect 66820 37508 66876 37510
rect 5800 34842 5856 34844
rect 5880 34842 5936 34844
rect 5960 34842 6016 34844
rect 6040 34842 6096 34844
rect 5800 34790 5846 34842
rect 5846 34790 5856 34842
rect 5880 34790 5910 34842
rect 5910 34790 5922 34842
rect 5922 34790 5936 34842
rect 5960 34790 5974 34842
rect 5974 34790 5986 34842
rect 5986 34790 6016 34842
rect 6040 34790 6050 34842
rect 6050 34790 6096 34842
rect 5800 34788 5856 34790
rect 5880 34788 5936 34790
rect 5960 34788 6016 34790
rect 6040 34788 6096 34790
rect 36520 34842 36576 34844
rect 36600 34842 36656 34844
rect 36680 34842 36736 34844
rect 36760 34842 36816 34844
rect 36520 34790 36566 34842
rect 36566 34790 36576 34842
rect 36600 34790 36630 34842
rect 36630 34790 36642 34842
rect 36642 34790 36656 34842
rect 36680 34790 36694 34842
rect 36694 34790 36706 34842
rect 36706 34790 36736 34842
rect 36760 34790 36770 34842
rect 36770 34790 36816 34842
rect 36520 34788 36576 34790
rect 36600 34788 36656 34790
rect 36680 34788 36736 34790
rect 36760 34788 36816 34790
rect 66580 36474 66636 36476
rect 66660 36474 66716 36476
rect 66740 36474 66796 36476
rect 66820 36474 66876 36476
rect 66580 36422 66626 36474
rect 66626 36422 66636 36474
rect 66660 36422 66690 36474
rect 66690 36422 66702 36474
rect 66702 36422 66716 36474
rect 66740 36422 66754 36474
rect 66754 36422 66766 36474
rect 66766 36422 66796 36474
rect 66820 36422 66830 36474
rect 66830 36422 66876 36474
rect 66580 36420 66636 36422
rect 66660 36420 66716 36422
rect 66740 36420 66796 36422
rect 66820 36420 66876 36422
rect 67240 39194 67296 39196
rect 67320 39194 67376 39196
rect 67400 39194 67456 39196
rect 67480 39194 67536 39196
rect 67240 39142 67286 39194
rect 67286 39142 67296 39194
rect 67320 39142 67350 39194
rect 67350 39142 67362 39194
rect 67362 39142 67376 39194
rect 67400 39142 67414 39194
rect 67414 39142 67426 39194
rect 67426 39142 67456 39194
rect 67480 39142 67490 39194
rect 67490 39142 67536 39194
rect 67240 39140 67296 39142
rect 67320 39140 67376 39142
rect 67400 39140 67456 39142
rect 67480 39140 67536 39142
rect 67240 38106 67296 38108
rect 67320 38106 67376 38108
rect 67400 38106 67456 38108
rect 67480 38106 67536 38108
rect 67240 38054 67286 38106
rect 67286 38054 67296 38106
rect 67320 38054 67350 38106
rect 67350 38054 67362 38106
rect 67362 38054 67376 38106
rect 67400 38054 67414 38106
rect 67414 38054 67426 38106
rect 67426 38054 67456 38106
rect 67480 38054 67490 38106
rect 67490 38054 67536 38106
rect 67240 38052 67296 38054
rect 67320 38052 67376 38054
rect 67400 38052 67456 38054
rect 67480 38052 67536 38054
rect 67240 37018 67296 37020
rect 67320 37018 67376 37020
rect 67400 37018 67456 37020
rect 67480 37018 67536 37020
rect 67240 36966 67286 37018
rect 67286 36966 67296 37018
rect 67320 36966 67350 37018
rect 67350 36966 67362 37018
rect 67362 36966 67376 37018
rect 67400 36966 67414 37018
rect 67414 36966 67426 37018
rect 67426 36966 67456 37018
rect 67480 36966 67490 37018
rect 67490 36966 67536 37018
rect 67240 36964 67296 36966
rect 67320 36964 67376 36966
rect 67400 36964 67456 36966
rect 67480 36964 67536 36966
rect 67240 35930 67296 35932
rect 67320 35930 67376 35932
rect 67400 35930 67456 35932
rect 67480 35930 67536 35932
rect 67240 35878 67286 35930
rect 67286 35878 67296 35930
rect 67320 35878 67350 35930
rect 67350 35878 67362 35930
rect 67362 35878 67376 35930
rect 67400 35878 67414 35930
rect 67414 35878 67426 35930
rect 67426 35878 67456 35930
rect 67480 35878 67490 35930
rect 67490 35878 67536 35930
rect 67240 35876 67296 35878
rect 67320 35876 67376 35878
rect 67400 35876 67456 35878
rect 67480 35876 67536 35878
rect 66580 35386 66636 35388
rect 66660 35386 66716 35388
rect 66740 35386 66796 35388
rect 66820 35386 66876 35388
rect 66580 35334 66626 35386
rect 66626 35334 66636 35386
rect 66660 35334 66690 35386
rect 66690 35334 66702 35386
rect 66702 35334 66716 35386
rect 66740 35334 66754 35386
rect 66754 35334 66766 35386
rect 66766 35334 66796 35386
rect 66820 35334 66830 35386
rect 66830 35334 66876 35386
rect 66580 35332 66636 35334
rect 66660 35332 66716 35334
rect 66740 35332 66796 35334
rect 66820 35332 66876 35334
rect 67240 34842 67296 34844
rect 67320 34842 67376 34844
rect 67400 34842 67456 34844
rect 67480 34842 67536 34844
rect 67240 34790 67286 34842
rect 67286 34790 67296 34842
rect 67320 34790 67350 34842
rect 67350 34790 67362 34842
rect 67362 34790 67376 34842
rect 67400 34790 67414 34842
rect 67414 34790 67426 34842
rect 67426 34790 67456 34842
rect 67480 34790 67490 34842
rect 67490 34790 67536 34842
rect 67240 34788 67296 34790
rect 67320 34788 67376 34790
rect 67400 34788 67456 34790
rect 67480 34788 67536 34790
rect 5140 34298 5196 34300
rect 5220 34298 5276 34300
rect 5300 34298 5356 34300
rect 5380 34298 5436 34300
rect 5140 34246 5186 34298
rect 5186 34246 5196 34298
rect 5220 34246 5250 34298
rect 5250 34246 5262 34298
rect 5262 34246 5276 34298
rect 5300 34246 5314 34298
rect 5314 34246 5326 34298
rect 5326 34246 5356 34298
rect 5380 34246 5390 34298
rect 5390 34246 5436 34298
rect 5140 34244 5196 34246
rect 5220 34244 5276 34246
rect 5300 34244 5356 34246
rect 5380 34244 5436 34246
rect 35860 34298 35916 34300
rect 35940 34298 35996 34300
rect 36020 34298 36076 34300
rect 36100 34298 36156 34300
rect 35860 34246 35906 34298
rect 35906 34246 35916 34298
rect 35940 34246 35970 34298
rect 35970 34246 35982 34298
rect 35982 34246 35996 34298
rect 36020 34246 36034 34298
rect 36034 34246 36046 34298
rect 36046 34246 36076 34298
rect 36100 34246 36110 34298
rect 36110 34246 36156 34298
rect 35860 34244 35916 34246
rect 35940 34244 35996 34246
rect 36020 34244 36076 34246
rect 36100 34244 36156 34246
rect 66580 34298 66636 34300
rect 66660 34298 66716 34300
rect 66740 34298 66796 34300
rect 66820 34298 66876 34300
rect 66580 34246 66626 34298
rect 66626 34246 66636 34298
rect 66660 34246 66690 34298
rect 66690 34246 66702 34298
rect 66702 34246 66716 34298
rect 66740 34246 66754 34298
rect 66754 34246 66766 34298
rect 66766 34246 66796 34298
rect 66820 34246 66830 34298
rect 66830 34246 66876 34298
rect 66580 34244 66636 34246
rect 66660 34244 66716 34246
rect 66740 34244 66796 34246
rect 66820 34244 66876 34246
rect 77482 38820 77538 38856
rect 77482 38800 77484 38820
rect 77484 38800 77536 38820
rect 77536 38800 77538 38820
rect 77482 38156 77484 38176
rect 77484 38156 77536 38176
rect 77536 38156 77538 38176
rect 77482 38120 77538 38156
rect 77482 37440 77538 37496
rect 77482 36760 77538 36816
rect 77482 34040 77538 34096
rect 5800 33754 5856 33756
rect 5880 33754 5936 33756
rect 5960 33754 6016 33756
rect 6040 33754 6096 33756
rect 5800 33702 5846 33754
rect 5846 33702 5856 33754
rect 5880 33702 5910 33754
rect 5910 33702 5922 33754
rect 5922 33702 5936 33754
rect 5960 33702 5974 33754
rect 5974 33702 5986 33754
rect 5986 33702 6016 33754
rect 6040 33702 6050 33754
rect 6050 33702 6096 33754
rect 5800 33700 5856 33702
rect 5880 33700 5936 33702
rect 5960 33700 6016 33702
rect 6040 33700 6096 33702
rect 36520 33754 36576 33756
rect 36600 33754 36656 33756
rect 36680 33754 36736 33756
rect 36760 33754 36816 33756
rect 36520 33702 36566 33754
rect 36566 33702 36576 33754
rect 36600 33702 36630 33754
rect 36630 33702 36642 33754
rect 36642 33702 36656 33754
rect 36680 33702 36694 33754
rect 36694 33702 36706 33754
rect 36706 33702 36736 33754
rect 36760 33702 36770 33754
rect 36770 33702 36816 33754
rect 36520 33700 36576 33702
rect 36600 33700 36656 33702
rect 36680 33700 36736 33702
rect 36760 33700 36816 33702
rect 67240 33754 67296 33756
rect 67320 33754 67376 33756
rect 67400 33754 67456 33756
rect 67480 33754 67536 33756
rect 67240 33702 67286 33754
rect 67286 33702 67296 33754
rect 67320 33702 67350 33754
rect 67350 33702 67362 33754
rect 67362 33702 67376 33754
rect 67400 33702 67414 33754
rect 67414 33702 67426 33754
rect 67426 33702 67456 33754
rect 67480 33702 67490 33754
rect 67490 33702 67536 33754
rect 67240 33700 67296 33702
rect 67320 33700 67376 33702
rect 67400 33700 67456 33702
rect 67480 33700 67536 33702
rect 5140 33210 5196 33212
rect 5220 33210 5276 33212
rect 5300 33210 5356 33212
rect 5380 33210 5436 33212
rect 5140 33158 5186 33210
rect 5186 33158 5196 33210
rect 5220 33158 5250 33210
rect 5250 33158 5262 33210
rect 5262 33158 5276 33210
rect 5300 33158 5314 33210
rect 5314 33158 5326 33210
rect 5326 33158 5356 33210
rect 5380 33158 5390 33210
rect 5390 33158 5436 33210
rect 5140 33156 5196 33158
rect 5220 33156 5276 33158
rect 5300 33156 5356 33158
rect 5380 33156 5436 33158
rect 35860 33210 35916 33212
rect 35940 33210 35996 33212
rect 36020 33210 36076 33212
rect 36100 33210 36156 33212
rect 35860 33158 35906 33210
rect 35906 33158 35916 33210
rect 35940 33158 35970 33210
rect 35970 33158 35982 33210
rect 35982 33158 35996 33210
rect 36020 33158 36034 33210
rect 36034 33158 36046 33210
rect 36046 33158 36076 33210
rect 36100 33158 36110 33210
rect 36110 33158 36156 33210
rect 35860 33156 35916 33158
rect 35940 33156 35996 33158
rect 36020 33156 36076 33158
rect 36100 33156 36156 33158
rect 66580 33210 66636 33212
rect 66660 33210 66716 33212
rect 66740 33210 66796 33212
rect 66820 33210 66876 33212
rect 66580 33158 66626 33210
rect 66626 33158 66636 33210
rect 66660 33158 66690 33210
rect 66690 33158 66702 33210
rect 66702 33158 66716 33210
rect 66740 33158 66754 33210
rect 66754 33158 66766 33210
rect 66766 33158 66796 33210
rect 66820 33158 66830 33210
rect 66830 33158 66876 33210
rect 66580 33156 66636 33158
rect 66660 33156 66716 33158
rect 66740 33156 66796 33158
rect 66820 33156 66876 33158
rect 5800 32666 5856 32668
rect 5880 32666 5936 32668
rect 5960 32666 6016 32668
rect 6040 32666 6096 32668
rect 5800 32614 5846 32666
rect 5846 32614 5856 32666
rect 5880 32614 5910 32666
rect 5910 32614 5922 32666
rect 5922 32614 5936 32666
rect 5960 32614 5974 32666
rect 5974 32614 5986 32666
rect 5986 32614 6016 32666
rect 6040 32614 6050 32666
rect 6050 32614 6096 32666
rect 5800 32612 5856 32614
rect 5880 32612 5936 32614
rect 5960 32612 6016 32614
rect 6040 32612 6096 32614
rect 36520 32666 36576 32668
rect 36600 32666 36656 32668
rect 36680 32666 36736 32668
rect 36760 32666 36816 32668
rect 36520 32614 36566 32666
rect 36566 32614 36576 32666
rect 36600 32614 36630 32666
rect 36630 32614 36642 32666
rect 36642 32614 36656 32666
rect 36680 32614 36694 32666
rect 36694 32614 36706 32666
rect 36706 32614 36736 32666
rect 36760 32614 36770 32666
rect 36770 32614 36816 32666
rect 36520 32612 36576 32614
rect 36600 32612 36656 32614
rect 36680 32612 36736 32614
rect 36760 32612 36816 32614
rect 67240 32666 67296 32668
rect 67320 32666 67376 32668
rect 67400 32666 67456 32668
rect 67480 32666 67536 32668
rect 67240 32614 67286 32666
rect 67286 32614 67296 32666
rect 67320 32614 67350 32666
rect 67350 32614 67362 32666
rect 67362 32614 67376 32666
rect 67400 32614 67414 32666
rect 67414 32614 67426 32666
rect 67426 32614 67456 32666
rect 67480 32614 67490 32666
rect 67490 32614 67536 32666
rect 67240 32612 67296 32614
rect 67320 32612 67376 32614
rect 67400 32612 67456 32614
rect 67480 32612 67536 32614
rect 5140 32122 5196 32124
rect 5220 32122 5276 32124
rect 5300 32122 5356 32124
rect 5380 32122 5436 32124
rect 5140 32070 5186 32122
rect 5186 32070 5196 32122
rect 5220 32070 5250 32122
rect 5250 32070 5262 32122
rect 5262 32070 5276 32122
rect 5300 32070 5314 32122
rect 5314 32070 5326 32122
rect 5326 32070 5356 32122
rect 5380 32070 5390 32122
rect 5390 32070 5436 32122
rect 5140 32068 5196 32070
rect 5220 32068 5276 32070
rect 5300 32068 5356 32070
rect 5380 32068 5436 32070
rect 35860 32122 35916 32124
rect 35940 32122 35996 32124
rect 36020 32122 36076 32124
rect 36100 32122 36156 32124
rect 35860 32070 35906 32122
rect 35906 32070 35916 32122
rect 35940 32070 35970 32122
rect 35970 32070 35982 32122
rect 35982 32070 35996 32122
rect 36020 32070 36034 32122
rect 36034 32070 36046 32122
rect 36046 32070 36076 32122
rect 36100 32070 36110 32122
rect 36110 32070 36156 32122
rect 35860 32068 35916 32070
rect 35940 32068 35996 32070
rect 36020 32068 36076 32070
rect 36100 32068 36156 32070
rect 66580 32122 66636 32124
rect 66660 32122 66716 32124
rect 66740 32122 66796 32124
rect 66820 32122 66876 32124
rect 66580 32070 66626 32122
rect 66626 32070 66636 32122
rect 66660 32070 66690 32122
rect 66690 32070 66702 32122
rect 66702 32070 66716 32122
rect 66740 32070 66754 32122
rect 66754 32070 66766 32122
rect 66766 32070 66796 32122
rect 66820 32070 66830 32122
rect 66830 32070 66876 32122
rect 66580 32068 66636 32070
rect 66660 32068 66716 32070
rect 66740 32068 66796 32070
rect 66820 32068 66876 32070
rect 1214 32000 1270 32056
rect 5800 31578 5856 31580
rect 5880 31578 5936 31580
rect 5960 31578 6016 31580
rect 6040 31578 6096 31580
rect 5800 31526 5846 31578
rect 5846 31526 5856 31578
rect 5880 31526 5910 31578
rect 5910 31526 5922 31578
rect 5922 31526 5936 31578
rect 5960 31526 5974 31578
rect 5974 31526 5986 31578
rect 5986 31526 6016 31578
rect 6040 31526 6050 31578
rect 6050 31526 6096 31578
rect 5800 31524 5856 31526
rect 5880 31524 5936 31526
rect 5960 31524 6016 31526
rect 6040 31524 6096 31526
rect 36520 31578 36576 31580
rect 36600 31578 36656 31580
rect 36680 31578 36736 31580
rect 36760 31578 36816 31580
rect 36520 31526 36566 31578
rect 36566 31526 36576 31578
rect 36600 31526 36630 31578
rect 36630 31526 36642 31578
rect 36642 31526 36656 31578
rect 36680 31526 36694 31578
rect 36694 31526 36706 31578
rect 36706 31526 36736 31578
rect 36760 31526 36770 31578
rect 36770 31526 36816 31578
rect 36520 31524 36576 31526
rect 36600 31524 36656 31526
rect 36680 31524 36736 31526
rect 36760 31524 36816 31526
rect 67240 31578 67296 31580
rect 67320 31578 67376 31580
rect 67400 31578 67456 31580
rect 67480 31578 67536 31580
rect 67240 31526 67286 31578
rect 67286 31526 67296 31578
rect 67320 31526 67350 31578
rect 67350 31526 67362 31578
rect 67362 31526 67376 31578
rect 67400 31526 67414 31578
rect 67414 31526 67426 31578
rect 67426 31526 67456 31578
rect 67480 31526 67490 31578
rect 67490 31526 67536 31578
rect 67240 31524 67296 31526
rect 67320 31524 67376 31526
rect 67400 31524 67456 31526
rect 67480 31524 67536 31526
rect 5140 31034 5196 31036
rect 5220 31034 5276 31036
rect 5300 31034 5356 31036
rect 5380 31034 5436 31036
rect 5140 30982 5186 31034
rect 5186 30982 5196 31034
rect 5220 30982 5250 31034
rect 5250 30982 5262 31034
rect 5262 30982 5276 31034
rect 5300 30982 5314 31034
rect 5314 30982 5326 31034
rect 5326 30982 5356 31034
rect 5380 30982 5390 31034
rect 5390 30982 5436 31034
rect 5140 30980 5196 30982
rect 5220 30980 5276 30982
rect 5300 30980 5356 30982
rect 5380 30980 5436 30982
rect 35860 31034 35916 31036
rect 35940 31034 35996 31036
rect 36020 31034 36076 31036
rect 36100 31034 36156 31036
rect 35860 30982 35906 31034
rect 35906 30982 35916 31034
rect 35940 30982 35970 31034
rect 35970 30982 35982 31034
rect 35982 30982 35996 31034
rect 36020 30982 36034 31034
rect 36034 30982 36046 31034
rect 36046 30982 36076 31034
rect 36100 30982 36110 31034
rect 36110 30982 36156 31034
rect 35860 30980 35916 30982
rect 35940 30980 35996 30982
rect 36020 30980 36076 30982
rect 36100 30980 36156 30982
rect 66580 31034 66636 31036
rect 66660 31034 66716 31036
rect 66740 31034 66796 31036
rect 66820 31034 66876 31036
rect 66580 30982 66626 31034
rect 66626 30982 66636 31034
rect 66660 30982 66690 31034
rect 66690 30982 66702 31034
rect 66702 30982 66716 31034
rect 66740 30982 66754 31034
rect 66754 30982 66766 31034
rect 66766 30982 66796 31034
rect 66820 30982 66830 31034
rect 66830 30982 66876 31034
rect 66580 30980 66636 30982
rect 66660 30980 66716 30982
rect 66740 30980 66796 30982
rect 66820 30980 66876 30982
rect 5800 30490 5856 30492
rect 5880 30490 5936 30492
rect 5960 30490 6016 30492
rect 6040 30490 6096 30492
rect 5800 30438 5846 30490
rect 5846 30438 5856 30490
rect 5880 30438 5910 30490
rect 5910 30438 5922 30490
rect 5922 30438 5936 30490
rect 5960 30438 5974 30490
rect 5974 30438 5986 30490
rect 5986 30438 6016 30490
rect 6040 30438 6050 30490
rect 6050 30438 6096 30490
rect 5800 30436 5856 30438
rect 5880 30436 5936 30438
rect 5960 30436 6016 30438
rect 6040 30436 6096 30438
rect 36520 30490 36576 30492
rect 36600 30490 36656 30492
rect 36680 30490 36736 30492
rect 36760 30490 36816 30492
rect 36520 30438 36566 30490
rect 36566 30438 36576 30490
rect 36600 30438 36630 30490
rect 36630 30438 36642 30490
rect 36642 30438 36656 30490
rect 36680 30438 36694 30490
rect 36694 30438 36706 30490
rect 36706 30438 36736 30490
rect 36760 30438 36770 30490
rect 36770 30438 36816 30490
rect 36520 30436 36576 30438
rect 36600 30436 36656 30438
rect 36680 30436 36736 30438
rect 36760 30436 36816 30438
rect 67240 30490 67296 30492
rect 67320 30490 67376 30492
rect 67400 30490 67456 30492
rect 67480 30490 67536 30492
rect 67240 30438 67286 30490
rect 67286 30438 67296 30490
rect 67320 30438 67350 30490
rect 67350 30438 67362 30490
rect 67362 30438 67376 30490
rect 67400 30438 67414 30490
rect 67414 30438 67426 30490
rect 67426 30438 67456 30490
rect 67480 30438 67490 30490
rect 67490 30438 67536 30490
rect 67240 30436 67296 30438
rect 67320 30436 67376 30438
rect 67400 30436 67456 30438
rect 67480 30436 67536 30438
rect 5140 29946 5196 29948
rect 5220 29946 5276 29948
rect 5300 29946 5356 29948
rect 5380 29946 5436 29948
rect 5140 29894 5186 29946
rect 5186 29894 5196 29946
rect 5220 29894 5250 29946
rect 5250 29894 5262 29946
rect 5262 29894 5276 29946
rect 5300 29894 5314 29946
rect 5314 29894 5326 29946
rect 5326 29894 5356 29946
rect 5380 29894 5390 29946
rect 5390 29894 5436 29946
rect 5140 29892 5196 29894
rect 5220 29892 5276 29894
rect 5300 29892 5356 29894
rect 5380 29892 5436 29894
rect 35860 29946 35916 29948
rect 35940 29946 35996 29948
rect 36020 29946 36076 29948
rect 36100 29946 36156 29948
rect 35860 29894 35906 29946
rect 35906 29894 35916 29946
rect 35940 29894 35970 29946
rect 35970 29894 35982 29946
rect 35982 29894 35996 29946
rect 36020 29894 36034 29946
rect 36034 29894 36046 29946
rect 36046 29894 36076 29946
rect 36100 29894 36110 29946
rect 36110 29894 36156 29946
rect 35860 29892 35916 29894
rect 35940 29892 35996 29894
rect 36020 29892 36076 29894
rect 36100 29892 36156 29894
rect 66580 29946 66636 29948
rect 66660 29946 66716 29948
rect 66740 29946 66796 29948
rect 66820 29946 66876 29948
rect 66580 29894 66626 29946
rect 66626 29894 66636 29946
rect 66660 29894 66690 29946
rect 66690 29894 66702 29946
rect 66702 29894 66716 29946
rect 66740 29894 66754 29946
rect 66754 29894 66766 29946
rect 66766 29894 66796 29946
rect 66820 29894 66830 29946
rect 66830 29894 66876 29946
rect 66580 29892 66636 29894
rect 66660 29892 66716 29894
rect 66740 29892 66796 29894
rect 66820 29892 66876 29894
rect 5800 29402 5856 29404
rect 5880 29402 5936 29404
rect 5960 29402 6016 29404
rect 6040 29402 6096 29404
rect 5800 29350 5846 29402
rect 5846 29350 5856 29402
rect 5880 29350 5910 29402
rect 5910 29350 5922 29402
rect 5922 29350 5936 29402
rect 5960 29350 5974 29402
rect 5974 29350 5986 29402
rect 5986 29350 6016 29402
rect 6040 29350 6050 29402
rect 6050 29350 6096 29402
rect 5800 29348 5856 29350
rect 5880 29348 5936 29350
rect 5960 29348 6016 29350
rect 6040 29348 6096 29350
rect 36520 29402 36576 29404
rect 36600 29402 36656 29404
rect 36680 29402 36736 29404
rect 36760 29402 36816 29404
rect 36520 29350 36566 29402
rect 36566 29350 36576 29402
rect 36600 29350 36630 29402
rect 36630 29350 36642 29402
rect 36642 29350 36656 29402
rect 36680 29350 36694 29402
rect 36694 29350 36706 29402
rect 36706 29350 36736 29402
rect 36760 29350 36770 29402
rect 36770 29350 36816 29402
rect 36520 29348 36576 29350
rect 36600 29348 36656 29350
rect 36680 29348 36736 29350
rect 36760 29348 36816 29350
rect 67240 29402 67296 29404
rect 67320 29402 67376 29404
rect 67400 29402 67456 29404
rect 67480 29402 67536 29404
rect 67240 29350 67286 29402
rect 67286 29350 67296 29402
rect 67320 29350 67350 29402
rect 67350 29350 67362 29402
rect 67362 29350 67376 29402
rect 67400 29350 67414 29402
rect 67414 29350 67426 29402
rect 67426 29350 67456 29402
rect 67480 29350 67490 29402
rect 67490 29350 67536 29402
rect 67240 29348 67296 29350
rect 67320 29348 67376 29350
rect 67400 29348 67456 29350
rect 67480 29348 67536 29350
rect 5140 28858 5196 28860
rect 5220 28858 5276 28860
rect 5300 28858 5356 28860
rect 5380 28858 5436 28860
rect 5140 28806 5186 28858
rect 5186 28806 5196 28858
rect 5220 28806 5250 28858
rect 5250 28806 5262 28858
rect 5262 28806 5276 28858
rect 5300 28806 5314 28858
rect 5314 28806 5326 28858
rect 5326 28806 5356 28858
rect 5380 28806 5390 28858
rect 5390 28806 5436 28858
rect 5140 28804 5196 28806
rect 5220 28804 5276 28806
rect 5300 28804 5356 28806
rect 5380 28804 5436 28806
rect 35860 28858 35916 28860
rect 35940 28858 35996 28860
rect 36020 28858 36076 28860
rect 36100 28858 36156 28860
rect 35860 28806 35906 28858
rect 35906 28806 35916 28858
rect 35940 28806 35970 28858
rect 35970 28806 35982 28858
rect 35982 28806 35996 28858
rect 36020 28806 36034 28858
rect 36034 28806 36046 28858
rect 36046 28806 36076 28858
rect 36100 28806 36110 28858
rect 36110 28806 36156 28858
rect 35860 28804 35916 28806
rect 35940 28804 35996 28806
rect 36020 28804 36076 28806
rect 36100 28804 36156 28806
rect 66580 28858 66636 28860
rect 66660 28858 66716 28860
rect 66740 28858 66796 28860
rect 66820 28858 66876 28860
rect 66580 28806 66626 28858
rect 66626 28806 66636 28858
rect 66660 28806 66690 28858
rect 66690 28806 66702 28858
rect 66702 28806 66716 28858
rect 66740 28806 66754 28858
rect 66754 28806 66766 28858
rect 66766 28806 66796 28858
rect 66820 28806 66830 28858
rect 66830 28806 66876 28858
rect 66580 28804 66636 28806
rect 66660 28804 66716 28806
rect 66740 28804 66796 28806
rect 66820 28804 66876 28806
rect 2318 28600 2374 28656
rect 5800 28314 5856 28316
rect 5880 28314 5936 28316
rect 5960 28314 6016 28316
rect 6040 28314 6096 28316
rect 5800 28262 5846 28314
rect 5846 28262 5856 28314
rect 5880 28262 5910 28314
rect 5910 28262 5922 28314
rect 5922 28262 5936 28314
rect 5960 28262 5974 28314
rect 5974 28262 5986 28314
rect 5986 28262 6016 28314
rect 6040 28262 6050 28314
rect 6050 28262 6096 28314
rect 5800 28260 5856 28262
rect 5880 28260 5936 28262
rect 5960 28260 6016 28262
rect 6040 28260 6096 28262
rect 36520 28314 36576 28316
rect 36600 28314 36656 28316
rect 36680 28314 36736 28316
rect 36760 28314 36816 28316
rect 36520 28262 36566 28314
rect 36566 28262 36576 28314
rect 36600 28262 36630 28314
rect 36630 28262 36642 28314
rect 36642 28262 36656 28314
rect 36680 28262 36694 28314
rect 36694 28262 36706 28314
rect 36706 28262 36736 28314
rect 36760 28262 36770 28314
rect 36770 28262 36816 28314
rect 36520 28260 36576 28262
rect 36600 28260 36656 28262
rect 36680 28260 36736 28262
rect 36760 28260 36816 28262
rect 67240 28314 67296 28316
rect 67320 28314 67376 28316
rect 67400 28314 67456 28316
rect 67480 28314 67536 28316
rect 67240 28262 67286 28314
rect 67286 28262 67296 28314
rect 67320 28262 67350 28314
rect 67350 28262 67362 28314
rect 67362 28262 67376 28314
rect 67400 28262 67414 28314
rect 67414 28262 67426 28314
rect 67426 28262 67456 28314
rect 67480 28262 67490 28314
rect 67490 28262 67536 28314
rect 67240 28260 67296 28262
rect 67320 28260 67376 28262
rect 67400 28260 67456 28262
rect 67480 28260 67536 28262
rect 1214 27956 1216 27976
rect 1216 27956 1268 27976
rect 1268 27956 1270 27976
rect 1214 27920 1270 27956
rect 5140 27770 5196 27772
rect 5220 27770 5276 27772
rect 5300 27770 5356 27772
rect 5380 27770 5436 27772
rect 5140 27718 5186 27770
rect 5186 27718 5196 27770
rect 5220 27718 5250 27770
rect 5250 27718 5262 27770
rect 5262 27718 5276 27770
rect 5300 27718 5314 27770
rect 5314 27718 5326 27770
rect 5326 27718 5356 27770
rect 5380 27718 5390 27770
rect 5390 27718 5436 27770
rect 5140 27716 5196 27718
rect 5220 27716 5276 27718
rect 5300 27716 5356 27718
rect 5380 27716 5436 27718
rect 35860 27770 35916 27772
rect 35940 27770 35996 27772
rect 36020 27770 36076 27772
rect 36100 27770 36156 27772
rect 35860 27718 35906 27770
rect 35906 27718 35916 27770
rect 35940 27718 35970 27770
rect 35970 27718 35982 27770
rect 35982 27718 35996 27770
rect 36020 27718 36034 27770
rect 36034 27718 36046 27770
rect 36046 27718 36076 27770
rect 36100 27718 36110 27770
rect 36110 27718 36156 27770
rect 35860 27716 35916 27718
rect 35940 27716 35996 27718
rect 36020 27716 36076 27718
rect 36100 27716 36156 27718
rect 66580 27770 66636 27772
rect 66660 27770 66716 27772
rect 66740 27770 66796 27772
rect 66820 27770 66876 27772
rect 66580 27718 66626 27770
rect 66626 27718 66636 27770
rect 66660 27718 66690 27770
rect 66690 27718 66702 27770
rect 66702 27718 66716 27770
rect 66740 27718 66754 27770
rect 66754 27718 66766 27770
rect 66766 27718 66796 27770
rect 66820 27718 66830 27770
rect 66830 27718 66876 27770
rect 66580 27716 66636 27718
rect 66660 27716 66716 27718
rect 66740 27716 66796 27718
rect 66820 27716 66876 27718
rect 5800 27226 5856 27228
rect 5880 27226 5936 27228
rect 5960 27226 6016 27228
rect 6040 27226 6096 27228
rect 5800 27174 5846 27226
rect 5846 27174 5856 27226
rect 5880 27174 5910 27226
rect 5910 27174 5922 27226
rect 5922 27174 5936 27226
rect 5960 27174 5974 27226
rect 5974 27174 5986 27226
rect 5986 27174 6016 27226
rect 6040 27174 6050 27226
rect 6050 27174 6096 27226
rect 5800 27172 5856 27174
rect 5880 27172 5936 27174
rect 5960 27172 6016 27174
rect 6040 27172 6096 27174
rect 36520 27226 36576 27228
rect 36600 27226 36656 27228
rect 36680 27226 36736 27228
rect 36760 27226 36816 27228
rect 36520 27174 36566 27226
rect 36566 27174 36576 27226
rect 36600 27174 36630 27226
rect 36630 27174 36642 27226
rect 36642 27174 36656 27226
rect 36680 27174 36694 27226
rect 36694 27174 36706 27226
rect 36706 27174 36736 27226
rect 36760 27174 36770 27226
rect 36770 27174 36816 27226
rect 36520 27172 36576 27174
rect 36600 27172 36656 27174
rect 36680 27172 36736 27174
rect 36760 27172 36816 27174
rect 67240 27226 67296 27228
rect 67320 27226 67376 27228
rect 67400 27226 67456 27228
rect 67480 27226 67536 27228
rect 67240 27174 67286 27226
rect 67286 27174 67296 27226
rect 67320 27174 67350 27226
rect 67350 27174 67362 27226
rect 67362 27174 67376 27226
rect 67400 27174 67414 27226
rect 67414 27174 67426 27226
rect 67426 27174 67456 27226
rect 67480 27174 67490 27226
rect 67490 27174 67536 27226
rect 67240 27172 67296 27174
rect 67320 27172 67376 27174
rect 67400 27172 67456 27174
rect 67480 27172 67536 27174
rect 5140 26682 5196 26684
rect 5220 26682 5276 26684
rect 5300 26682 5356 26684
rect 5380 26682 5436 26684
rect 5140 26630 5186 26682
rect 5186 26630 5196 26682
rect 5220 26630 5250 26682
rect 5250 26630 5262 26682
rect 5262 26630 5276 26682
rect 5300 26630 5314 26682
rect 5314 26630 5326 26682
rect 5326 26630 5356 26682
rect 5380 26630 5390 26682
rect 5390 26630 5436 26682
rect 5140 26628 5196 26630
rect 5220 26628 5276 26630
rect 5300 26628 5356 26630
rect 5380 26628 5436 26630
rect 35860 26682 35916 26684
rect 35940 26682 35996 26684
rect 36020 26682 36076 26684
rect 36100 26682 36156 26684
rect 35860 26630 35906 26682
rect 35906 26630 35916 26682
rect 35940 26630 35970 26682
rect 35970 26630 35982 26682
rect 35982 26630 35996 26682
rect 36020 26630 36034 26682
rect 36034 26630 36046 26682
rect 36046 26630 36076 26682
rect 36100 26630 36110 26682
rect 36110 26630 36156 26682
rect 35860 26628 35916 26630
rect 35940 26628 35996 26630
rect 36020 26628 36076 26630
rect 36100 26628 36156 26630
rect 66580 26682 66636 26684
rect 66660 26682 66716 26684
rect 66740 26682 66796 26684
rect 66820 26682 66876 26684
rect 66580 26630 66626 26682
rect 66626 26630 66636 26682
rect 66660 26630 66690 26682
rect 66690 26630 66702 26682
rect 66702 26630 66716 26682
rect 66740 26630 66754 26682
rect 66754 26630 66766 26682
rect 66766 26630 66796 26682
rect 66820 26630 66830 26682
rect 66830 26630 66876 26682
rect 66580 26628 66636 26630
rect 66660 26628 66716 26630
rect 66740 26628 66796 26630
rect 66820 26628 66876 26630
rect 1214 26560 1270 26616
rect 5800 26138 5856 26140
rect 5880 26138 5936 26140
rect 5960 26138 6016 26140
rect 6040 26138 6096 26140
rect 5800 26086 5846 26138
rect 5846 26086 5856 26138
rect 5880 26086 5910 26138
rect 5910 26086 5922 26138
rect 5922 26086 5936 26138
rect 5960 26086 5974 26138
rect 5974 26086 5986 26138
rect 5986 26086 6016 26138
rect 6040 26086 6050 26138
rect 6050 26086 6096 26138
rect 5800 26084 5856 26086
rect 5880 26084 5936 26086
rect 5960 26084 6016 26086
rect 6040 26084 6096 26086
rect 36520 26138 36576 26140
rect 36600 26138 36656 26140
rect 36680 26138 36736 26140
rect 36760 26138 36816 26140
rect 36520 26086 36566 26138
rect 36566 26086 36576 26138
rect 36600 26086 36630 26138
rect 36630 26086 36642 26138
rect 36642 26086 36656 26138
rect 36680 26086 36694 26138
rect 36694 26086 36706 26138
rect 36706 26086 36736 26138
rect 36760 26086 36770 26138
rect 36770 26086 36816 26138
rect 36520 26084 36576 26086
rect 36600 26084 36656 26086
rect 36680 26084 36736 26086
rect 36760 26084 36816 26086
rect 67240 26138 67296 26140
rect 67320 26138 67376 26140
rect 67400 26138 67456 26140
rect 67480 26138 67536 26140
rect 67240 26086 67286 26138
rect 67286 26086 67296 26138
rect 67320 26086 67350 26138
rect 67350 26086 67362 26138
rect 67362 26086 67376 26138
rect 67400 26086 67414 26138
rect 67414 26086 67426 26138
rect 67426 26086 67456 26138
rect 67480 26086 67490 26138
rect 67490 26086 67536 26138
rect 67240 26084 67296 26086
rect 67320 26084 67376 26086
rect 67400 26084 67456 26086
rect 67480 26084 67536 26086
rect 2318 25880 2374 25936
rect 5140 25594 5196 25596
rect 5220 25594 5276 25596
rect 5300 25594 5356 25596
rect 5380 25594 5436 25596
rect 5140 25542 5186 25594
rect 5186 25542 5196 25594
rect 5220 25542 5250 25594
rect 5250 25542 5262 25594
rect 5262 25542 5276 25594
rect 5300 25542 5314 25594
rect 5314 25542 5326 25594
rect 5326 25542 5356 25594
rect 5380 25542 5390 25594
rect 5390 25542 5436 25594
rect 5140 25540 5196 25542
rect 5220 25540 5276 25542
rect 5300 25540 5356 25542
rect 5380 25540 5436 25542
rect 35860 25594 35916 25596
rect 35940 25594 35996 25596
rect 36020 25594 36076 25596
rect 36100 25594 36156 25596
rect 35860 25542 35906 25594
rect 35906 25542 35916 25594
rect 35940 25542 35970 25594
rect 35970 25542 35982 25594
rect 35982 25542 35996 25594
rect 36020 25542 36034 25594
rect 36034 25542 36046 25594
rect 36046 25542 36076 25594
rect 36100 25542 36110 25594
rect 36110 25542 36156 25594
rect 35860 25540 35916 25542
rect 35940 25540 35996 25542
rect 36020 25540 36076 25542
rect 36100 25540 36156 25542
rect 66580 25594 66636 25596
rect 66660 25594 66716 25596
rect 66740 25594 66796 25596
rect 66820 25594 66876 25596
rect 66580 25542 66626 25594
rect 66626 25542 66636 25594
rect 66660 25542 66690 25594
rect 66690 25542 66702 25594
rect 66702 25542 66716 25594
rect 66740 25542 66754 25594
rect 66754 25542 66766 25594
rect 66766 25542 66796 25594
rect 66820 25542 66830 25594
rect 66830 25542 66876 25594
rect 66580 25540 66636 25542
rect 66660 25540 66716 25542
rect 66740 25540 66796 25542
rect 66820 25540 66876 25542
rect 5800 25050 5856 25052
rect 5880 25050 5936 25052
rect 5960 25050 6016 25052
rect 6040 25050 6096 25052
rect 5800 24998 5846 25050
rect 5846 24998 5856 25050
rect 5880 24998 5910 25050
rect 5910 24998 5922 25050
rect 5922 24998 5936 25050
rect 5960 24998 5974 25050
rect 5974 24998 5986 25050
rect 5986 24998 6016 25050
rect 6040 24998 6050 25050
rect 6050 24998 6096 25050
rect 5800 24996 5856 24998
rect 5880 24996 5936 24998
rect 5960 24996 6016 24998
rect 6040 24996 6096 24998
rect 36520 25050 36576 25052
rect 36600 25050 36656 25052
rect 36680 25050 36736 25052
rect 36760 25050 36816 25052
rect 36520 24998 36566 25050
rect 36566 24998 36576 25050
rect 36600 24998 36630 25050
rect 36630 24998 36642 25050
rect 36642 24998 36656 25050
rect 36680 24998 36694 25050
rect 36694 24998 36706 25050
rect 36706 24998 36736 25050
rect 36760 24998 36770 25050
rect 36770 24998 36816 25050
rect 36520 24996 36576 24998
rect 36600 24996 36656 24998
rect 36680 24996 36736 24998
rect 36760 24996 36816 24998
rect 67240 25050 67296 25052
rect 67320 25050 67376 25052
rect 67400 25050 67456 25052
rect 67480 25050 67536 25052
rect 67240 24998 67286 25050
rect 67286 24998 67296 25050
rect 67320 24998 67350 25050
rect 67350 24998 67362 25050
rect 67362 24998 67376 25050
rect 67400 24998 67414 25050
rect 67414 24998 67426 25050
rect 67426 24998 67456 25050
rect 67480 24998 67490 25050
rect 67490 24998 67536 25050
rect 67240 24996 67296 24998
rect 67320 24996 67376 24998
rect 67400 24996 67456 24998
rect 67480 24996 67536 24998
rect 5140 24506 5196 24508
rect 5220 24506 5276 24508
rect 5300 24506 5356 24508
rect 5380 24506 5436 24508
rect 5140 24454 5186 24506
rect 5186 24454 5196 24506
rect 5220 24454 5250 24506
rect 5250 24454 5262 24506
rect 5262 24454 5276 24506
rect 5300 24454 5314 24506
rect 5314 24454 5326 24506
rect 5326 24454 5356 24506
rect 5380 24454 5390 24506
rect 5390 24454 5436 24506
rect 5140 24452 5196 24454
rect 5220 24452 5276 24454
rect 5300 24452 5356 24454
rect 5380 24452 5436 24454
rect 35860 24506 35916 24508
rect 35940 24506 35996 24508
rect 36020 24506 36076 24508
rect 36100 24506 36156 24508
rect 35860 24454 35906 24506
rect 35906 24454 35916 24506
rect 35940 24454 35970 24506
rect 35970 24454 35982 24506
rect 35982 24454 35996 24506
rect 36020 24454 36034 24506
rect 36034 24454 36046 24506
rect 36046 24454 36076 24506
rect 36100 24454 36110 24506
rect 36110 24454 36156 24506
rect 35860 24452 35916 24454
rect 35940 24452 35996 24454
rect 36020 24452 36076 24454
rect 36100 24452 36156 24454
rect 66580 24506 66636 24508
rect 66660 24506 66716 24508
rect 66740 24506 66796 24508
rect 66820 24506 66876 24508
rect 66580 24454 66626 24506
rect 66626 24454 66636 24506
rect 66660 24454 66690 24506
rect 66690 24454 66702 24506
rect 66702 24454 66716 24506
rect 66740 24454 66754 24506
rect 66754 24454 66766 24506
rect 66766 24454 66796 24506
rect 66820 24454 66830 24506
rect 66830 24454 66876 24506
rect 66580 24452 66636 24454
rect 66660 24452 66716 24454
rect 66740 24452 66796 24454
rect 66820 24452 66876 24454
rect 5800 23962 5856 23964
rect 5880 23962 5936 23964
rect 5960 23962 6016 23964
rect 6040 23962 6096 23964
rect 5800 23910 5846 23962
rect 5846 23910 5856 23962
rect 5880 23910 5910 23962
rect 5910 23910 5922 23962
rect 5922 23910 5936 23962
rect 5960 23910 5974 23962
rect 5974 23910 5986 23962
rect 5986 23910 6016 23962
rect 6040 23910 6050 23962
rect 6050 23910 6096 23962
rect 5800 23908 5856 23910
rect 5880 23908 5936 23910
rect 5960 23908 6016 23910
rect 6040 23908 6096 23910
rect 36520 23962 36576 23964
rect 36600 23962 36656 23964
rect 36680 23962 36736 23964
rect 36760 23962 36816 23964
rect 36520 23910 36566 23962
rect 36566 23910 36576 23962
rect 36600 23910 36630 23962
rect 36630 23910 36642 23962
rect 36642 23910 36656 23962
rect 36680 23910 36694 23962
rect 36694 23910 36706 23962
rect 36706 23910 36736 23962
rect 36760 23910 36770 23962
rect 36770 23910 36816 23962
rect 36520 23908 36576 23910
rect 36600 23908 36656 23910
rect 36680 23908 36736 23910
rect 36760 23908 36816 23910
rect 67240 23962 67296 23964
rect 67320 23962 67376 23964
rect 67400 23962 67456 23964
rect 67480 23962 67536 23964
rect 67240 23910 67286 23962
rect 67286 23910 67296 23962
rect 67320 23910 67350 23962
rect 67350 23910 67362 23962
rect 67362 23910 67376 23962
rect 67400 23910 67414 23962
rect 67414 23910 67426 23962
rect 67426 23910 67456 23962
rect 67480 23910 67490 23962
rect 67490 23910 67536 23962
rect 67240 23908 67296 23910
rect 67320 23908 67376 23910
rect 67400 23908 67456 23910
rect 67480 23908 67536 23910
rect 5140 23418 5196 23420
rect 5220 23418 5276 23420
rect 5300 23418 5356 23420
rect 5380 23418 5436 23420
rect 5140 23366 5186 23418
rect 5186 23366 5196 23418
rect 5220 23366 5250 23418
rect 5250 23366 5262 23418
rect 5262 23366 5276 23418
rect 5300 23366 5314 23418
rect 5314 23366 5326 23418
rect 5326 23366 5356 23418
rect 5380 23366 5390 23418
rect 5390 23366 5436 23418
rect 5140 23364 5196 23366
rect 5220 23364 5276 23366
rect 5300 23364 5356 23366
rect 5380 23364 5436 23366
rect 35860 23418 35916 23420
rect 35940 23418 35996 23420
rect 36020 23418 36076 23420
rect 36100 23418 36156 23420
rect 35860 23366 35906 23418
rect 35906 23366 35916 23418
rect 35940 23366 35970 23418
rect 35970 23366 35982 23418
rect 35982 23366 35996 23418
rect 36020 23366 36034 23418
rect 36034 23366 36046 23418
rect 36046 23366 36076 23418
rect 36100 23366 36110 23418
rect 36110 23366 36156 23418
rect 35860 23364 35916 23366
rect 35940 23364 35996 23366
rect 36020 23364 36076 23366
rect 36100 23364 36156 23366
rect 66580 23418 66636 23420
rect 66660 23418 66716 23420
rect 66740 23418 66796 23420
rect 66820 23418 66876 23420
rect 66580 23366 66626 23418
rect 66626 23366 66636 23418
rect 66660 23366 66690 23418
rect 66690 23366 66702 23418
rect 66702 23366 66716 23418
rect 66740 23366 66754 23418
rect 66754 23366 66766 23418
rect 66766 23366 66796 23418
rect 66820 23366 66830 23418
rect 66830 23366 66876 23418
rect 66580 23364 66636 23366
rect 66660 23364 66716 23366
rect 66740 23364 66796 23366
rect 66820 23364 66876 23366
rect 2318 23160 2374 23216
rect 5800 22874 5856 22876
rect 5880 22874 5936 22876
rect 5960 22874 6016 22876
rect 6040 22874 6096 22876
rect 5800 22822 5846 22874
rect 5846 22822 5856 22874
rect 5880 22822 5910 22874
rect 5910 22822 5922 22874
rect 5922 22822 5936 22874
rect 5960 22822 5974 22874
rect 5974 22822 5986 22874
rect 5986 22822 6016 22874
rect 6040 22822 6050 22874
rect 6050 22822 6096 22874
rect 5800 22820 5856 22822
rect 5880 22820 5936 22822
rect 5960 22820 6016 22822
rect 6040 22820 6096 22822
rect 36520 22874 36576 22876
rect 36600 22874 36656 22876
rect 36680 22874 36736 22876
rect 36760 22874 36816 22876
rect 36520 22822 36566 22874
rect 36566 22822 36576 22874
rect 36600 22822 36630 22874
rect 36630 22822 36642 22874
rect 36642 22822 36656 22874
rect 36680 22822 36694 22874
rect 36694 22822 36706 22874
rect 36706 22822 36736 22874
rect 36760 22822 36770 22874
rect 36770 22822 36816 22874
rect 36520 22820 36576 22822
rect 36600 22820 36656 22822
rect 36680 22820 36736 22822
rect 36760 22820 36816 22822
rect 67240 22874 67296 22876
rect 67320 22874 67376 22876
rect 67400 22874 67456 22876
rect 67480 22874 67536 22876
rect 67240 22822 67286 22874
rect 67286 22822 67296 22874
rect 67320 22822 67350 22874
rect 67350 22822 67362 22874
rect 67362 22822 67376 22874
rect 67400 22822 67414 22874
rect 67414 22822 67426 22874
rect 67426 22822 67456 22874
rect 67480 22822 67490 22874
rect 67490 22822 67536 22874
rect 67240 22820 67296 22822
rect 67320 22820 67376 22822
rect 67400 22820 67456 22822
rect 67480 22820 67536 22822
rect 5140 22330 5196 22332
rect 5220 22330 5276 22332
rect 5300 22330 5356 22332
rect 5380 22330 5436 22332
rect 5140 22278 5186 22330
rect 5186 22278 5196 22330
rect 5220 22278 5250 22330
rect 5250 22278 5262 22330
rect 5262 22278 5276 22330
rect 5300 22278 5314 22330
rect 5314 22278 5326 22330
rect 5326 22278 5356 22330
rect 5380 22278 5390 22330
rect 5390 22278 5436 22330
rect 5140 22276 5196 22278
rect 5220 22276 5276 22278
rect 5300 22276 5356 22278
rect 5380 22276 5436 22278
rect 35860 22330 35916 22332
rect 35940 22330 35996 22332
rect 36020 22330 36076 22332
rect 36100 22330 36156 22332
rect 35860 22278 35906 22330
rect 35906 22278 35916 22330
rect 35940 22278 35970 22330
rect 35970 22278 35982 22330
rect 35982 22278 35996 22330
rect 36020 22278 36034 22330
rect 36034 22278 36046 22330
rect 36046 22278 36076 22330
rect 36100 22278 36110 22330
rect 36110 22278 36156 22330
rect 35860 22276 35916 22278
rect 35940 22276 35996 22278
rect 36020 22276 36076 22278
rect 36100 22276 36156 22278
rect 66580 22330 66636 22332
rect 66660 22330 66716 22332
rect 66740 22330 66796 22332
rect 66820 22330 66876 22332
rect 66580 22278 66626 22330
rect 66626 22278 66636 22330
rect 66660 22278 66690 22330
rect 66690 22278 66702 22330
rect 66702 22278 66716 22330
rect 66740 22278 66754 22330
rect 66754 22278 66766 22330
rect 66766 22278 66796 22330
rect 66820 22278 66830 22330
rect 66830 22278 66876 22330
rect 66580 22276 66636 22278
rect 66660 22276 66716 22278
rect 66740 22276 66796 22278
rect 66820 22276 66876 22278
rect 5800 21786 5856 21788
rect 5880 21786 5936 21788
rect 5960 21786 6016 21788
rect 6040 21786 6096 21788
rect 5800 21734 5846 21786
rect 5846 21734 5856 21786
rect 5880 21734 5910 21786
rect 5910 21734 5922 21786
rect 5922 21734 5936 21786
rect 5960 21734 5974 21786
rect 5974 21734 5986 21786
rect 5986 21734 6016 21786
rect 6040 21734 6050 21786
rect 6050 21734 6096 21786
rect 5800 21732 5856 21734
rect 5880 21732 5936 21734
rect 5960 21732 6016 21734
rect 6040 21732 6096 21734
rect 36520 21786 36576 21788
rect 36600 21786 36656 21788
rect 36680 21786 36736 21788
rect 36760 21786 36816 21788
rect 36520 21734 36566 21786
rect 36566 21734 36576 21786
rect 36600 21734 36630 21786
rect 36630 21734 36642 21786
rect 36642 21734 36656 21786
rect 36680 21734 36694 21786
rect 36694 21734 36706 21786
rect 36706 21734 36736 21786
rect 36760 21734 36770 21786
rect 36770 21734 36816 21786
rect 36520 21732 36576 21734
rect 36600 21732 36656 21734
rect 36680 21732 36736 21734
rect 36760 21732 36816 21734
rect 67240 21786 67296 21788
rect 67320 21786 67376 21788
rect 67400 21786 67456 21788
rect 67480 21786 67536 21788
rect 67240 21734 67286 21786
rect 67286 21734 67296 21786
rect 67320 21734 67350 21786
rect 67350 21734 67362 21786
rect 67362 21734 67376 21786
rect 67400 21734 67414 21786
rect 67414 21734 67426 21786
rect 67426 21734 67456 21786
rect 67480 21734 67490 21786
rect 67490 21734 67536 21786
rect 67240 21732 67296 21734
rect 67320 21732 67376 21734
rect 67400 21732 67456 21734
rect 67480 21732 67536 21734
rect 5140 21242 5196 21244
rect 5220 21242 5276 21244
rect 5300 21242 5356 21244
rect 5380 21242 5436 21244
rect 5140 21190 5186 21242
rect 5186 21190 5196 21242
rect 5220 21190 5250 21242
rect 5250 21190 5262 21242
rect 5262 21190 5276 21242
rect 5300 21190 5314 21242
rect 5314 21190 5326 21242
rect 5326 21190 5356 21242
rect 5380 21190 5390 21242
rect 5390 21190 5436 21242
rect 5140 21188 5196 21190
rect 5220 21188 5276 21190
rect 5300 21188 5356 21190
rect 5380 21188 5436 21190
rect 35860 21242 35916 21244
rect 35940 21242 35996 21244
rect 36020 21242 36076 21244
rect 36100 21242 36156 21244
rect 35860 21190 35906 21242
rect 35906 21190 35916 21242
rect 35940 21190 35970 21242
rect 35970 21190 35982 21242
rect 35982 21190 35996 21242
rect 36020 21190 36034 21242
rect 36034 21190 36046 21242
rect 36046 21190 36076 21242
rect 36100 21190 36110 21242
rect 36110 21190 36156 21242
rect 35860 21188 35916 21190
rect 35940 21188 35996 21190
rect 36020 21188 36076 21190
rect 36100 21188 36156 21190
rect 66580 21242 66636 21244
rect 66660 21242 66716 21244
rect 66740 21242 66796 21244
rect 66820 21242 66876 21244
rect 66580 21190 66626 21242
rect 66626 21190 66636 21242
rect 66660 21190 66690 21242
rect 66690 21190 66702 21242
rect 66702 21190 66716 21242
rect 66740 21190 66754 21242
rect 66754 21190 66766 21242
rect 66766 21190 66796 21242
rect 66820 21190 66830 21242
rect 66830 21190 66876 21242
rect 66580 21188 66636 21190
rect 66660 21188 66716 21190
rect 66740 21188 66796 21190
rect 66820 21188 66876 21190
rect 77574 21120 77630 21176
rect 5800 20698 5856 20700
rect 5880 20698 5936 20700
rect 5960 20698 6016 20700
rect 6040 20698 6096 20700
rect 5800 20646 5846 20698
rect 5846 20646 5856 20698
rect 5880 20646 5910 20698
rect 5910 20646 5922 20698
rect 5922 20646 5936 20698
rect 5960 20646 5974 20698
rect 5974 20646 5986 20698
rect 5986 20646 6016 20698
rect 6040 20646 6050 20698
rect 6050 20646 6096 20698
rect 5800 20644 5856 20646
rect 5880 20644 5936 20646
rect 5960 20644 6016 20646
rect 6040 20644 6096 20646
rect 36520 20698 36576 20700
rect 36600 20698 36656 20700
rect 36680 20698 36736 20700
rect 36760 20698 36816 20700
rect 36520 20646 36566 20698
rect 36566 20646 36576 20698
rect 36600 20646 36630 20698
rect 36630 20646 36642 20698
rect 36642 20646 36656 20698
rect 36680 20646 36694 20698
rect 36694 20646 36706 20698
rect 36706 20646 36736 20698
rect 36760 20646 36770 20698
rect 36770 20646 36816 20698
rect 36520 20644 36576 20646
rect 36600 20644 36656 20646
rect 36680 20644 36736 20646
rect 36760 20644 36816 20646
rect 67240 20698 67296 20700
rect 67320 20698 67376 20700
rect 67400 20698 67456 20700
rect 67480 20698 67536 20700
rect 67240 20646 67286 20698
rect 67286 20646 67296 20698
rect 67320 20646 67350 20698
rect 67350 20646 67362 20698
rect 67362 20646 67376 20698
rect 67400 20646 67414 20698
rect 67414 20646 67426 20698
rect 67426 20646 67456 20698
rect 67480 20646 67490 20698
rect 67490 20646 67536 20698
rect 67240 20644 67296 20646
rect 67320 20644 67376 20646
rect 67400 20644 67456 20646
rect 67480 20644 67536 20646
rect 5140 20154 5196 20156
rect 5220 20154 5276 20156
rect 5300 20154 5356 20156
rect 5380 20154 5436 20156
rect 5140 20102 5186 20154
rect 5186 20102 5196 20154
rect 5220 20102 5250 20154
rect 5250 20102 5262 20154
rect 5262 20102 5276 20154
rect 5300 20102 5314 20154
rect 5314 20102 5326 20154
rect 5326 20102 5356 20154
rect 5380 20102 5390 20154
rect 5390 20102 5436 20154
rect 5140 20100 5196 20102
rect 5220 20100 5276 20102
rect 5300 20100 5356 20102
rect 5380 20100 5436 20102
rect 35860 20154 35916 20156
rect 35940 20154 35996 20156
rect 36020 20154 36076 20156
rect 36100 20154 36156 20156
rect 35860 20102 35906 20154
rect 35906 20102 35916 20154
rect 35940 20102 35970 20154
rect 35970 20102 35982 20154
rect 35982 20102 35996 20154
rect 36020 20102 36034 20154
rect 36034 20102 36046 20154
rect 36046 20102 36076 20154
rect 36100 20102 36110 20154
rect 36110 20102 36156 20154
rect 35860 20100 35916 20102
rect 35940 20100 35996 20102
rect 36020 20100 36076 20102
rect 36100 20100 36156 20102
rect 66580 20154 66636 20156
rect 66660 20154 66716 20156
rect 66740 20154 66796 20156
rect 66820 20154 66876 20156
rect 66580 20102 66626 20154
rect 66626 20102 66636 20154
rect 66660 20102 66690 20154
rect 66690 20102 66702 20154
rect 66702 20102 66716 20154
rect 66740 20102 66754 20154
rect 66754 20102 66766 20154
rect 66766 20102 66796 20154
rect 66820 20102 66830 20154
rect 66830 20102 66876 20154
rect 66580 20100 66636 20102
rect 66660 20100 66716 20102
rect 66740 20100 66796 20102
rect 66820 20100 66876 20102
rect 5800 19610 5856 19612
rect 5880 19610 5936 19612
rect 5960 19610 6016 19612
rect 6040 19610 6096 19612
rect 5800 19558 5846 19610
rect 5846 19558 5856 19610
rect 5880 19558 5910 19610
rect 5910 19558 5922 19610
rect 5922 19558 5936 19610
rect 5960 19558 5974 19610
rect 5974 19558 5986 19610
rect 5986 19558 6016 19610
rect 6040 19558 6050 19610
rect 6050 19558 6096 19610
rect 5800 19556 5856 19558
rect 5880 19556 5936 19558
rect 5960 19556 6016 19558
rect 6040 19556 6096 19558
rect 36520 19610 36576 19612
rect 36600 19610 36656 19612
rect 36680 19610 36736 19612
rect 36760 19610 36816 19612
rect 36520 19558 36566 19610
rect 36566 19558 36576 19610
rect 36600 19558 36630 19610
rect 36630 19558 36642 19610
rect 36642 19558 36656 19610
rect 36680 19558 36694 19610
rect 36694 19558 36706 19610
rect 36706 19558 36736 19610
rect 36760 19558 36770 19610
rect 36770 19558 36816 19610
rect 36520 19556 36576 19558
rect 36600 19556 36656 19558
rect 36680 19556 36736 19558
rect 36760 19556 36816 19558
rect 67240 19610 67296 19612
rect 67320 19610 67376 19612
rect 67400 19610 67456 19612
rect 67480 19610 67536 19612
rect 67240 19558 67286 19610
rect 67286 19558 67296 19610
rect 67320 19558 67350 19610
rect 67350 19558 67362 19610
rect 67362 19558 67376 19610
rect 67400 19558 67414 19610
rect 67414 19558 67426 19610
rect 67426 19558 67456 19610
rect 67480 19558 67490 19610
rect 67490 19558 67536 19610
rect 67240 19556 67296 19558
rect 67320 19556 67376 19558
rect 67400 19556 67456 19558
rect 67480 19556 67536 19558
rect 5140 19066 5196 19068
rect 5220 19066 5276 19068
rect 5300 19066 5356 19068
rect 5380 19066 5436 19068
rect 5140 19014 5186 19066
rect 5186 19014 5196 19066
rect 5220 19014 5250 19066
rect 5250 19014 5262 19066
rect 5262 19014 5276 19066
rect 5300 19014 5314 19066
rect 5314 19014 5326 19066
rect 5326 19014 5356 19066
rect 5380 19014 5390 19066
rect 5390 19014 5436 19066
rect 5140 19012 5196 19014
rect 5220 19012 5276 19014
rect 5300 19012 5356 19014
rect 5380 19012 5436 19014
rect 35860 19066 35916 19068
rect 35940 19066 35996 19068
rect 36020 19066 36076 19068
rect 36100 19066 36156 19068
rect 35860 19014 35906 19066
rect 35906 19014 35916 19066
rect 35940 19014 35970 19066
rect 35970 19014 35982 19066
rect 35982 19014 35996 19066
rect 36020 19014 36034 19066
rect 36034 19014 36046 19066
rect 36046 19014 36076 19066
rect 36100 19014 36110 19066
rect 36110 19014 36156 19066
rect 35860 19012 35916 19014
rect 35940 19012 35996 19014
rect 36020 19012 36076 19014
rect 36100 19012 36156 19014
rect 66580 19066 66636 19068
rect 66660 19066 66716 19068
rect 66740 19066 66796 19068
rect 66820 19066 66876 19068
rect 66580 19014 66626 19066
rect 66626 19014 66636 19066
rect 66660 19014 66690 19066
rect 66690 19014 66702 19066
rect 66702 19014 66716 19066
rect 66740 19014 66754 19066
rect 66754 19014 66766 19066
rect 66766 19014 66796 19066
rect 66820 19014 66830 19066
rect 66830 19014 66876 19066
rect 66580 19012 66636 19014
rect 66660 19012 66716 19014
rect 66740 19012 66796 19014
rect 66820 19012 66876 19014
rect 5800 18522 5856 18524
rect 5880 18522 5936 18524
rect 5960 18522 6016 18524
rect 6040 18522 6096 18524
rect 5800 18470 5846 18522
rect 5846 18470 5856 18522
rect 5880 18470 5910 18522
rect 5910 18470 5922 18522
rect 5922 18470 5936 18522
rect 5960 18470 5974 18522
rect 5974 18470 5986 18522
rect 5986 18470 6016 18522
rect 6040 18470 6050 18522
rect 6050 18470 6096 18522
rect 5800 18468 5856 18470
rect 5880 18468 5936 18470
rect 5960 18468 6016 18470
rect 6040 18468 6096 18470
rect 36520 18522 36576 18524
rect 36600 18522 36656 18524
rect 36680 18522 36736 18524
rect 36760 18522 36816 18524
rect 36520 18470 36566 18522
rect 36566 18470 36576 18522
rect 36600 18470 36630 18522
rect 36630 18470 36642 18522
rect 36642 18470 36656 18522
rect 36680 18470 36694 18522
rect 36694 18470 36706 18522
rect 36706 18470 36736 18522
rect 36760 18470 36770 18522
rect 36770 18470 36816 18522
rect 36520 18468 36576 18470
rect 36600 18468 36656 18470
rect 36680 18468 36736 18470
rect 36760 18468 36816 18470
rect 67240 18522 67296 18524
rect 67320 18522 67376 18524
rect 67400 18522 67456 18524
rect 67480 18522 67536 18524
rect 67240 18470 67286 18522
rect 67286 18470 67296 18522
rect 67320 18470 67350 18522
rect 67350 18470 67362 18522
rect 67362 18470 67376 18522
rect 67400 18470 67414 18522
rect 67414 18470 67426 18522
rect 67426 18470 67456 18522
rect 67480 18470 67490 18522
rect 67490 18470 67536 18522
rect 67240 18468 67296 18470
rect 67320 18468 67376 18470
rect 67400 18468 67456 18470
rect 67480 18468 67536 18470
rect 5140 17978 5196 17980
rect 5220 17978 5276 17980
rect 5300 17978 5356 17980
rect 5380 17978 5436 17980
rect 5140 17926 5186 17978
rect 5186 17926 5196 17978
rect 5220 17926 5250 17978
rect 5250 17926 5262 17978
rect 5262 17926 5276 17978
rect 5300 17926 5314 17978
rect 5314 17926 5326 17978
rect 5326 17926 5356 17978
rect 5380 17926 5390 17978
rect 5390 17926 5436 17978
rect 5140 17924 5196 17926
rect 5220 17924 5276 17926
rect 5300 17924 5356 17926
rect 5380 17924 5436 17926
rect 35860 17978 35916 17980
rect 35940 17978 35996 17980
rect 36020 17978 36076 17980
rect 36100 17978 36156 17980
rect 35860 17926 35906 17978
rect 35906 17926 35916 17978
rect 35940 17926 35970 17978
rect 35970 17926 35982 17978
rect 35982 17926 35996 17978
rect 36020 17926 36034 17978
rect 36034 17926 36046 17978
rect 36046 17926 36076 17978
rect 36100 17926 36110 17978
rect 36110 17926 36156 17978
rect 35860 17924 35916 17926
rect 35940 17924 35996 17926
rect 36020 17924 36076 17926
rect 36100 17924 36156 17926
rect 66580 17978 66636 17980
rect 66660 17978 66716 17980
rect 66740 17978 66796 17980
rect 66820 17978 66876 17980
rect 66580 17926 66626 17978
rect 66626 17926 66636 17978
rect 66660 17926 66690 17978
rect 66690 17926 66702 17978
rect 66702 17926 66716 17978
rect 66740 17926 66754 17978
rect 66754 17926 66766 17978
rect 66766 17926 66796 17978
rect 66820 17926 66830 17978
rect 66830 17926 66876 17978
rect 66580 17924 66636 17926
rect 66660 17924 66716 17926
rect 66740 17924 66796 17926
rect 66820 17924 66876 17926
rect 5800 17434 5856 17436
rect 5880 17434 5936 17436
rect 5960 17434 6016 17436
rect 6040 17434 6096 17436
rect 5800 17382 5846 17434
rect 5846 17382 5856 17434
rect 5880 17382 5910 17434
rect 5910 17382 5922 17434
rect 5922 17382 5936 17434
rect 5960 17382 5974 17434
rect 5974 17382 5986 17434
rect 5986 17382 6016 17434
rect 6040 17382 6050 17434
rect 6050 17382 6096 17434
rect 5800 17380 5856 17382
rect 5880 17380 5936 17382
rect 5960 17380 6016 17382
rect 6040 17380 6096 17382
rect 36520 17434 36576 17436
rect 36600 17434 36656 17436
rect 36680 17434 36736 17436
rect 36760 17434 36816 17436
rect 36520 17382 36566 17434
rect 36566 17382 36576 17434
rect 36600 17382 36630 17434
rect 36630 17382 36642 17434
rect 36642 17382 36656 17434
rect 36680 17382 36694 17434
rect 36694 17382 36706 17434
rect 36706 17382 36736 17434
rect 36760 17382 36770 17434
rect 36770 17382 36816 17434
rect 36520 17380 36576 17382
rect 36600 17380 36656 17382
rect 36680 17380 36736 17382
rect 36760 17380 36816 17382
rect 67240 17434 67296 17436
rect 67320 17434 67376 17436
rect 67400 17434 67456 17436
rect 67480 17434 67536 17436
rect 67240 17382 67286 17434
rect 67286 17382 67296 17434
rect 67320 17382 67350 17434
rect 67350 17382 67362 17434
rect 67362 17382 67376 17434
rect 67400 17382 67414 17434
rect 67414 17382 67426 17434
rect 67426 17382 67456 17434
rect 67480 17382 67490 17434
rect 67490 17382 67536 17434
rect 67240 17380 67296 17382
rect 67320 17380 67376 17382
rect 67400 17380 67456 17382
rect 67480 17380 67536 17382
rect 5140 16890 5196 16892
rect 5220 16890 5276 16892
rect 5300 16890 5356 16892
rect 5380 16890 5436 16892
rect 5140 16838 5186 16890
rect 5186 16838 5196 16890
rect 5220 16838 5250 16890
rect 5250 16838 5262 16890
rect 5262 16838 5276 16890
rect 5300 16838 5314 16890
rect 5314 16838 5326 16890
rect 5326 16838 5356 16890
rect 5380 16838 5390 16890
rect 5390 16838 5436 16890
rect 5140 16836 5196 16838
rect 5220 16836 5276 16838
rect 5300 16836 5356 16838
rect 5380 16836 5436 16838
rect 35860 16890 35916 16892
rect 35940 16890 35996 16892
rect 36020 16890 36076 16892
rect 36100 16890 36156 16892
rect 35860 16838 35906 16890
rect 35906 16838 35916 16890
rect 35940 16838 35970 16890
rect 35970 16838 35982 16890
rect 35982 16838 35996 16890
rect 36020 16838 36034 16890
rect 36034 16838 36046 16890
rect 36046 16838 36076 16890
rect 36100 16838 36110 16890
rect 36110 16838 36156 16890
rect 35860 16836 35916 16838
rect 35940 16836 35996 16838
rect 36020 16836 36076 16838
rect 36100 16836 36156 16838
rect 66580 16890 66636 16892
rect 66660 16890 66716 16892
rect 66740 16890 66796 16892
rect 66820 16890 66876 16892
rect 66580 16838 66626 16890
rect 66626 16838 66636 16890
rect 66660 16838 66690 16890
rect 66690 16838 66702 16890
rect 66702 16838 66716 16890
rect 66740 16838 66754 16890
rect 66754 16838 66766 16890
rect 66766 16838 66796 16890
rect 66820 16838 66830 16890
rect 66830 16838 66876 16890
rect 66580 16836 66636 16838
rect 66660 16836 66716 16838
rect 66740 16836 66796 16838
rect 66820 16836 66876 16838
rect 77574 16360 77630 16416
rect 5800 16346 5856 16348
rect 5880 16346 5936 16348
rect 5960 16346 6016 16348
rect 6040 16346 6096 16348
rect 5800 16294 5846 16346
rect 5846 16294 5856 16346
rect 5880 16294 5910 16346
rect 5910 16294 5922 16346
rect 5922 16294 5936 16346
rect 5960 16294 5974 16346
rect 5974 16294 5986 16346
rect 5986 16294 6016 16346
rect 6040 16294 6050 16346
rect 6050 16294 6096 16346
rect 5800 16292 5856 16294
rect 5880 16292 5936 16294
rect 5960 16292 6016 16294
rect 6040 16292 6096 16294
rect 36520 16346 36576 16348
rect 36600 16346 36656 16348
rect 36680 16346 36736 16348
rect 36760 16346 36816 16348
rect 36520 16294 36566 16346
rect 36566 16294 36576 16346
rect 36600 16294 36630 16346
rect 36630 16294 36642 16346
rect 36642 16294 36656 16346
rect 36680 16294 36694 16346
rect 36694 16294 36706 16346
rect 36706 16294 36736 16346
rect 36760 16294 36770 16346
rect 36770 16294 36816 16346
rect 36520 16292 36576 16294
rect 36600 16292 36656 16294
rect 36680 16292 36736 16294
rect 36760 16292 36816 16294
rect 67240 16346 67296 16348
rect 67320 16346 67376 16348
rect 67400 16346 67456 16348
rect 67480 16346 67536 16348
rect 67240 16294 67286 16346
rect 67286 16294 67296 16346
rect 67320 16294 67350 16346
rect 67350 16294 67362 16346
rect 67362 16294 67376 16346
rect 67400 16294 67414 16346
rect 67414 16294 67426 16346
rect 67426 16294 67456 16346
rect 67480 16294 67490 16346
rect 67490 16294 67536 16346
rect 67240 16292 67296 16294
rect 67320 16292 67376 16294
rect 67400 16292 67456 16294
rect 67480 16292 67536 16294
rect 5140 15802 5196 15804
rect 5220 15802 5276 15804
rect 5300 15802 5356 15804
rect 5380 15802 5436 15804
rect 5140 15750 5186 15802
rect 5186 15750 5196 15802
rect 5220 15750 5250 15802
rect 5250 15750 5262 15802
rect 5262 15750 5276 15802
rect 5300 15750 5314 15802
rect 5314 15750 5326 15802
rect 5326 15750 5356 15802
rect 5380 15750 5390 15802
rect 5390 15750 5436 15802
rect 5140 15748 5196 15750
rect 5220 15748 5276 15750
rect 5300 15748 5356 15750
rect 5380 15748 5436 15750
rect 35860 15802 35916 15804
rect 35940 15802 35996 15804
rect 36020 15802 36076 15804
rect 36100 15802 36156 15804
rect 35860 15750 35906 15802
rect 35906 15750 35916 15802
rect 35940 15750 35970 15802
rect 35970 15750 35982 15802
rect 35982 15750 35996 15802
rect 36020 15750 36034 15802
rect 36034 15750 36046 15802
rect 36046 15750 36076 15802
rect 36100 15750 36110 15802
rect 36110 15750 36156 15802
rect 35860 15748 35916 15750
rect 35940 15748 35996 15750
rect 36020 15748 36076 15750
rect 36100 15748 36156 15750
rect 66580 15802 66636 15804
rect 66660 15802 66716 15804
rect 66740 15802 66796 15804
rect 66820 15802 66876 15804
rect 66580 15750 66626 15802
rect 66626 15750 66636 15802
rect 66660 15750 66690 15802
rect 66690 15750 66702 15802
rect 66702 15750 66716 15802
rect 66740 15750 66754 15802
rect 66754 15750 66766 15802
rect 66766 15750 66796 15802
rect 66820 15750 66830 15802
rect 66830 15750 66876 15802
rect 66580 15748 66636 15750
rect 66660 15748 66716 15750
rect 66740 15748 66796 15750
rect 66820 15748 66876 15750
rect 5800 15258 5856 15260
rect 5880 15258 5936 15260
rect 5960 15258 6016 15260
rect 6040 15258 6096 15260
rect 5800 15206 5846 15258
rect 5846 15206 5856 15258
rect 5880 15206 5910 15258
rect 5910 15206 5922 15258
rect 5922 15206 5936 15258
rect 5960 15206 5974 15258
rect 5974 15206 5986 15258
rect 5986 15206 6016 15258
rect 6040 15206 6050 15258
rect 6050 15206 6096 15258
rect 5800 15204 5856 15206
rect 5880 15204 5936 15206
rect 5960 15204 6016 15206
rect 6040 15204 6096 15206
rect 36520 15258 36576 15260
rect 36600 15258 36656 15260
rect 36680 15258 36736 15260
rect 36760 15258 36816 15260
rect 36520 15206 36566 15258
rect 36566 15206 36576 15258
rect 36600 15206 36630 15258
rect 36630 15206 36642 15258
rect 36642 15206 36656 15258
rect 36680 15206 36694 15258
rect 36694 15206 36706 15258
rect 36706 15206 36736 15258
rect 36760 15206 36770 15258
rect 36770 15206 36816 15258
rect 36520 15204 36576 15206
rect 36600 15204 36656 15206
rect 36680 15204 36736 15206
rect 36760 15204 36816 15206
rect 67240 15258 67296 15260
rect 67320 15258 67376 15260
rect 67400 15258 67456 15260
rect 67480 15258 67536 15260
rect 67240 15206 67286 15258
rect 67286 15206 67296 15258
rect 67320 15206 67350 15258
rect 67350 15206 67362 15258
rect 67362 15206 67376 15258
rect 67400 15206 67414 15258
rect 67414 15206 67426 15258
rect 67426 15206 67456 15258
rect 67480 15206 67490 15258
rect 67490 15206 67536 15258
rect 67240 15204 67296 15206
rect 67320 15204 67376 15206
rect 67400 15204 67456 15206
rect 67480 15204 67536 15206
rect 5140 14714 5196 14716
rect 5220 14714 5276 14716
rect 5300 14714 5356 14716
rect 5380 14714 5436 14716
rect 5140 14662 5186 14714
rect 5186 14662 5196 14714
rect 5220 14662 5250 14714
rect 5250 14662 5262 14714
rect 5262 14662 5276 14714
rect 5300 14662 5314 14714
rect 5314 14662 5326 14714
rect 5326 14662 5356 14714
rect 5380 14662 5390 14714
rect 5390 14662 5436 14714
rect 5140 14660 5196 14662
rect 5220 14660 5276 14662
rect 5300 14660 5356 14662
rect 5380 14660 5436 14662
rect 35860 14714 35916 14716
rect 35940 14714 35996 14716
rect 36020 14714 36076 14716
rect 36100 14714 36156 14716
rect 35860 14662 35906 14714
rect 35906 14662 35916 14714
rect 35940 14662 35970 14714
rect 35970 14662 35982 14714
rect 35982 14662 35996 14714
rect 36020 14662 36034 14714
rect 36034 14662 36046 14714
rect 36046 14662 36076 14714
rect 36100 14662 36110 14714
rect 36110 14662 36156 14714
rect 35860 14660 35916 14662
rect 35940 14660 35996 14662
rect 36020 14660 36076 14662
rect 36100 14660 36156 14662
rect 66580 14714 66636 14716
rect 66660 14714 66716 14716
rect 66740 14714 66796 14716
rect 66820 14714 66876 14716
rect 66580 14662 66626 14714
rect 66626 14662 66636 14714
rect 66660 14662 66690 14714
rect 66690 14662 66702 14714
rect 66702 14662 66716 14714
rect 66740 14662 66754 14714
rect 66754 14662 66766 14714
rect 66766 14662 66796 14714
rect 66820 14662 66830 14714
rect 66830 14662 66876 14714
rect 66580 14660 66636 14662
rect 66660 14660 66716 14662
rect 66740 14660 66796 14662
rect 66820 14660 66876 14662
rect 5800 14170 5856 14172
rect 5880 14170 5936 14172
rect 5960 14170 6016 14172
rect 6040 14170 6096 14172
rect 5800 14118 5846 14170
rect 5846 14118 5856 14170
rect 5880 14118 5910 14170
rect 5910 14118 5922 14170
rect 5922 14118 5936 14170
rect 5960 14118 5974 14170
rect 5974 14118 5986 14170
rect 5986 14118 6016 14170
rect 6040 14118 6050 14170
rect 6050 14118 6096 14170
rect 5800 14116 5856 14118
rect 5880 14116 5936 14118
rect 5960 14116 6016 14118
rect 6040 14116 6096 14118
rect 36520 14170 36576 14172
rect 36600 14170 36656 14172
rect 36680 14170 36736 14172
rect 36760 14170 36816 14172
rect 36520 14118 36566 14170
rect 36566 14118 36576 14170
rect 36600 14118 36630 14170
rect 36630 14118 36642 14170
rect 36642 14118 36656 14170
rect 36680 14118 36694 14170
rect 36694 14118 36706 14170
rect 36706 14118 36736 14170
rect 36760 14118 36770 14170
rect 36770 14118 36816 14170
rect 36520 14116 36576 14118
rect 36600 14116 36656 14118
rect 36680 14116 36736 14118
rect 36760 14116 36816 14118
rect 67240 14170 67296 14172
rect 67320 14170 67376 14172
rect 67400 14170 67456 14172
rect 67480 14170 67536 14172
rect 67240 14118 67286 14170
rect 67286 14118 67296 14170
rect 67320 14118 67350 14170
rect 67350 14118 67362 14170
rect 67362 14118 67376 14170
rect 67400 14118 67414 14170
rect 67414 14118 67426 14170
rect 67426 14118 67456 14170
rect 67480 14118 67490 14170
rect 67490 14118 67536 14170
rect 67240 14116 67296 14118
rect 67320 14116 67376 14118
rect 67400 14116 67456 14118
rect 67480 14116 67536 14118
rect 5140 13626 5196 13628
rect 5220 13626 5276 13628
rect 5300 13626 5356 13628
rect 5380 13626 5436 13628
rect 5140 13574 5186 13626
rect 5186 13574 5196 13626
rect 5220 13574 5250 13626
rect 5250 13574 5262 13626
rect 5262 13574 5276 13626
rect 5300 13574 5314 13626
rect 5314 13574 5326 13626
rect 5326 13574 5356 13626
rect 5380 13574 5390 13626
rect 5390 13574 5436 13626
rect 5140 13572 5196 13574
rect 5220 13572 5276 13574
rect 5300 13572 5356 13574
rect 5380 13572 5436 13574
rect 35860 13626 35916 13628
rect 35940 13626 35996 13628
rect 36020 13626 36076 13628
rect 36100 13626 36156 13628
rect 35860 13574 35906 13626
rect 35906 13574 35916 13626
rect 35940 13574 35970 13626
rect 35970 13574 35982 13626
rect 35982 13574 35996 13626
rect 36020 13574 36034 13626
rect 36034 13574 36046 13626
rect 36046 13574 36076 13626
rect 36100 13574 36110 13626
rect 36110 13574 36156 13626
rect 35860 13572 35916 13574
rect 35940 13572 35996 13574
rect 36020 13572 36076 13574
rect 36100 13572 36156 13574
rect 66580 13626 66636 13628
rect 66660 13626 66716 13628
rect 66740 13626 66796 13628
rect 66820 13626 66876 13628
rect 66580 13574 66626 13626
rect 66626 13574 66636 13626
rect 66660 13574 66690 13626
rect 66690 13574 66702 13626
rect 66702 13574 66716 13626
rect 66740 13574 66754 13626
rect 66754 13574 66766 13626
rect 66766 13574 66796 13626
rect 66820 13574 66830 13626
rect 66830 13574 66876 13626
rect 66580 13572 66636 13574
rect 66660 13572 66716 13574
rect 66740 13572 66796 13574
rect 66820 13572 66876 13574
rect 5800 13082 5856 13084
rect 5880 13082 5936 13084
rect 5960 13082 6016 13084
rect 6040 13082 6096 13084
rect 5800 13030 5846 13082
rect 5846 13030 5856 13082
rect 5880 13030 5910 13082
rect 5910 13030 5922 13082
rect 5922 13030 5936 13082
rect 5960 13030 5974 13082
rect 5974 13030 5986 13082
rect 5986 13030 6016 13082
rect 6040 13030 6050 13082
rect 6050 13030 6096 13082
rect 5800 13028 5856 13030
rect 5880 13028 5936 13030
rect 5960 13028 6016 13030
rect 6040 13028 6096 13030
rect 36520 13082 36576 13084
rect 36600 13082 36656 13084
rect 36680 13082 36736 13084
rect 36760 13082 36816 13084
rect 36520 13030 36566 13082
rect 36566 13030 36576 13082
rect 36600 13030 36630 13082
rect 36630 13030 36642 13082
rect 36642 13030 36656 13082
rect 36680 13030 36694 13082
rect 36694 13030 36706 13082
rect 36706 13030 36736 13082
rect 36760 13030 36770 13082
rect 36770 13030 36816 13082
rect 36520 13028 36576 13030
rect 36600 13028 36656 13030
rect 36680 13028 36736 13030
rect 36760 13028 36816 13030
rect 67240 13082 67296 13084
rect 67320 13082 67376 13084
rect 67400 13082 67456 13084
rect 67480 13082 67536 13084
rect 67240 13030 67286 13082
rect 67286 13030 67296 13082
rect 67320 13030 67350 13082
rect 67350 13030 67362 13082
rect 67362 13030 67376 13082
rect 67400 13030 67414 13082
rect 67414 13030 67426 13082
rect 67426 13030 67456 13082
rect 67480 13030 67490 13082
rect 67490 13030 67536 13082
rect 67240 13028 67296 13030
rect 67320 13028 67376 13030
rect 67400 13028 67456 13030
rect 67480 13028 67536 13030
rect 5140 12538 5196 12540
rect 5220 12538 5276 12540
rect 5300 12538 5356 12540
rect 5380 12538 5436 12540
rect 5140 12486 5186 12538
rect 5186 12486 5196 12538
rect 5220 12486 5250 12538
rect 5250 12486 5262 12538
rect 5262 12486 5276 12538
rect 5300 12486 5314 12538
rect 5314 12486 5326 12538
rect 5326 12486 5356 12538
rect 5380 12486 5390 12538
rect 5390 12486 5436 12538
rect 5140 12484 5196 12486
rect 5220 12484 5276 12486
rect 5300 12484 5356 12486
rect 5380 12484 5436 12486
rect 35860 12538 35916 12540
rect 35940 12538 35996 12540
rect 36020 12538 36076 12540
rect 36100 12538 36156 12540
rect 35860 12486 35906 12538
rect 35906 12486 35916 12538
rect 35940 12486 35970 12538
rect 35970 12486 35982 12538
rect 35982 12486 35996 12538
rect 36020 12486 36034 12538
rect 36034 12486 36046 12538
rect 36046 12486 36076 12538
rect 36100 12486 36110 12538
rect 36110 12486 36156 12538
rect 35860 12484 35916 12486
rect 35940 12484 35996 12486
rect 36020 12484 36076 12486
rect 36100 12484 36156 12486
rect 66580 12538 66636 12540
rect 66660 12538 66716 12540
rect 66740 12538 66796 12540
rect 66820 12538 66876 12540
rect 66580 12486 66626 12538
rect 66626 12486 66636 12538
rect 66660 12486 66690 12538
rect 66690 12486 66702 12538
rect 66702 12486 66716 12538
rect 66740 12486 66754 12538
rect 66754 12486 66766 12538
rect 66766 12486 66796 12538
rect 66820 12486 66830 12538
rect 66830 12486 66876 12538
rect 66580 12484 66636 12486
rect 66660 12484 66716 12486
rect 66740 12484 66796 12486
rect 66820 12484 66876 12486
rect 5800 11994 5856 11996
rect 5880 11994 5936 11996
rect 5960 11994 6016 11996
rect 6040 11994 6096 11996
rect 5800 11942 5846 11994
rect 5846 11942 5856 11994
rect 5880 11942 5910 11994
rect 5910 11942 5922 11994
rect 5922 11942 5936 11994
rect 5960 11942 5974 11994
rect 5974 11942 5986 11994
rect 5986 11942 6016 11994
rect 6040 11942 6050 11994
rect 6050 11942 6096 11994
rect 5800 11940 5856 11942
rect 5880 11940 5936 11942
rect 5960 11940 6016 11942
rect 6040 11940 6096 11942
rect 36520 11994 36576 11996
rect 36600 11994 36656 11996
rect 36680 11994 36736 11996
rect 36760 11994 36816 11996
rect 36520 11942 36566 11994
rect 36566 11942 36576 11994
rect 36600 11942 36630 11994
rect 36630 11942 36642 11994
rect 36642 11942 36656 11994
rect 36680 11942 36694 11994
rect 36694 11942 36706 11994
rect 36706 11942 36736 11994
rect 36760 11942 36770 11994
rect 36770 11942 36816 11994
rect 36520 11940 36576 11942
rect 36600 11940 36656 11942
rect 36680 11940 36736 11942
rect 36760 11940 36816 11942
rect 67240 11994 67296 11996
rect 67320 11994 67376 11996
rect 67400 11994 67456 11996
rect 67480 11994 67536 11996
rect 67240 11942 67286 11994
rect 67286 11942 67296 11994
rect 67320 11942 67350 11994
rect 67350 11942 67362 11994
rect 67362 11942 67376 11994
rect 67400 11942 67414 11994
rect 67414 11942 67426 11994
rect 67426 11942 67456 11994
rect 67480 11942 67490 11994
rect 67490 11942 67536 11994
rect 67240 11940 67296 11942
rect 67320 11940 67376 11942
rect 67400 11940 67456 11942
rect 67480 11940 67536 11942
rect 5140 11450 5196 11452
rect 5220 11450 5276 11452
rect 5300 11450 5356 11452
rect 5380 11450 5436 11452
rect 5140 11398 5186 11450
rect 5186 11398 5196 11450
rect 5220 11398 5250 11450
rect 5250 11398 5262 11450
rect 5262 11398 5276 11450
rect 5300 11398 5314 11450
rect 5314 11398 5326 11450
rect 5326 11398 5356 11450
rect 5380 11398 5390 11450
rect 5390 11398 5436 11450
rect 5140 11396 5196 11398
rect 5220 11396 5276 11398
rect 5300 11396 5356 11398
rect 5380 11396 5436 11398
rect 35860 11450 35916 11452
rect 35940 11450 35996 11452
rect 36020 11450 36076 11452
rect 36100 11450 36156 11452
rect 35860 11398 35906 11450
rect 35906 11398 35916 11450
rect 35940 11398 35970 11450
rect 35970 11398 35982 11450
rect 35982 11398 35996 11450
rect 36020 11398 36034 11450
rect 36034 11398 36046 11450
rect 36046 11398 36076 11450
rect 36100 11398 36110 11450
rect 36110 11398 36156 11450
rect 35860 11396 35916 11398
rect 35940 11396 35996 11398
rect 36020 11396 36076 11398
rect 36100 11396 36156 11398
rect 66580 11450 66636 11452
rect 66660 11450 66716 11452
rect 66740 11450 66796 11452
rect 66820 11450 66876 11452
rect 66580 11398 66626 11450
rect 66626 11398 66636 11450
rect 66660 11398 66690 11450
rect 66690 11398 66702 11450
rect 66702 11398 66716 11450
rect 66740 11398 66754 11450
rect 66754 11398 66766 11450
rect 66766 11398 66796 11450
rect 66820 11398 66830 11450
rect 66830 11398 66876 11450
rect 66580 11396 66636 11398
rect 66660 11396 66716 11398
rect 66740 11396 66796 11398
rect 66820 11396 66876 11398
rect 5800 10906 5856 10908
rect 5880 10906 5936 10908
rect 5960 10906 6016 10908
rect 6040 10906 6096 10908
rect 5800 10854 5846 10906
rect 5846 10854 5856 10906
rect 5880 10854 5910 10906
rect 5910 10854 5922 10906
rect 5922 10854 5936 10906
rect 5960 10854 5974 10906
rect 5974 10854 5986 10906
rect 5986 10854 6016 10906
rect 6040 10854 6050 10906
rect 6050 10854 6096 10906
rect 5800 10852 5856 10854
rect 5880 10852 5936 10854
rect 5960 10852 6016 10854
rect 6040 10852 6096 10854
rect 36520 10906 36576 10908
rect 36600 10906 36656 10908
rect 36680 10906 36736 10908
rect 36760 10906 36816 10908
rect 36520 10854 36566 10906
rect 36566 10854 36576 10906
rect 36600 10854 36630 10906
rect 36630 10854 36642 10906
rect 36642 10854 36656 10906
rect 36680 10854 36694 10906
rect 36694 10854 36706 10906
rect 36706 10854 36736 10906
rect 36760 10854 36770 10906
rect 36770 10854 36816 10906
rect 36520 10852 36576 10854
rect 36600 10852 36656 10854
rect 36680 10852 36736 10854
rect 36760 10852 36816 10854
rect 67240 10906 67296 10908
rect 67320 10906 67376 10908
rect 67400 10906 67456 10908
rect 67480 10906 67536 10908
rect 67240 10854 67286 10906
rect 67286 10854 67296 10906
rect 67320 10854 67350 10906
rect 67350 10854 67362 10906
rect 67362 10854 67376 10906
rect 67400 10854 67414 10906
rect 67414 10854 67426 10906
rect 67426 10854 67456 10906
rect 67480 10854 67490 10906
rect 67490 10854 67536 10906
rect 67240 10852 67296 10854
rect 67320 10852 67376 10854
rect 67400 10852 67456 10854
rect 67480 10852 67536 10854
rect 5140 10362 5196 10364
rect 5220 10362 5276 10364
rect 5300 10362 5356 10364
rect 5380 10362 5436 10364
rect 5140 10310 5186 10362
rect 5186 10310 5196 10362
rect 5220 10310 5250 10362
rect 5250 10310 5262 10362
rect 5262 10310 5276 10362
rect 5300 10310 5314 10362
rect 5314 10310 5326 10362
rect 5326 10310 5356 10362
rect 5380 10310 5390 10362
rect 5390 10310 5436 10362
rect 5140 10308 5196 10310
rect 5220 10308 5276 10310
rect 5300 10308 5356 10310
rect 5380 10308 5436 10310
rect 35860 10362 35916 10364
rect 35940 10362 35996 10364
rect 36020 10362 36076 10364
rect 36100 10362 36156 10364
rect 35860 10310 35906 10362
rect 35906 10310 35916 10362
rect 35940 10310 35970 10362
rect 35970 10310 35982 10362
rect 35982 10310 35996 10362
rect 36020 10310 36034 10362
rect 36034 10310 36046 10362
rect 36046 10310 36076 10362
rect 36100 10310 36110 10362
rect 36110 10310 36156 10362
rect 35860 10308 35916 10310
rect 35940 10308 35996 10310
rect 36020 10308 36076 10310
rect 36100 10308 36156 10310
rect 66580 10362 66636 10364
rect 66660 10362 66716 10364
rect 66740 10362 66796 10364
rect 66820 10362 66876 10364
rect 66580 10310 66626 10362
rect 66626 10310 66636 10362
rect 66660 10310 66690 10362
rect 66690 10310 66702 10362
rect 66702 10310 66716 10362
rect 66740 10310 66754 10362
rect 66754 10310 66766 10362
rect 66766 10310 66796 10362
rect 66820 10310 66830 10362
rect 66830 10310 66876 10362
rect 66580 10308 66636 10310
rect 66660 10308 66716 10310
rect 66740 10308 66796 10310
rect 66820 10308 66876 10310
rect 5800 9818 5856 9820
rect 5880 9818 5936 9820
rect 5960 9818 6016 9820
rect 6040 9818 6096 9820
rect 5800 9766 5846 9818
rect 5846 9766 5856 9818
rect 5880 9766 5910 9818
rect 5910 9766 5922 9818
rect 5922 9766 5936 9818
rect 5960 9766 5974 9818
rect 5974 9766 5986 9818
rect 5986 9766 6016 9818
rect 6040 9766 6050 9818
rect 6050 9766 6096 9818
rect 5800 9764 5856 9766
rect 5880 9764 5936 9766
rect 5960 9764 6016 9766
rect 6040 9764 6096 9766
rect 36520 9818 36576 9820
rect 36600 9818 36656 9820
rect 36680 9818 36736 9820
rect 36760 9818 36816 9820
rect 36520 9766 36566 9818
rect 36566 9766 36576 9818
rect 36600 9766 36630 9818
rect 36630 9766 36642 9818
rect 36642 9766 36656 9818
rect 36680 9766 36694 9818
rect 36694 9766 36706 9818
rect 36706 9766 36736 9818
rect 36760 9766 36770 9818
rect 36770 9766 36816 9818
rect 36520 9764 36576 9766
rect 36600 9764 36656 9766
rect 36680 9764 36736 9766
rect 36760 9764 36816 9766
rect 67240 9818 67296 9820
rect 67320 9818 67376 9820
rect 67400 9818 67456 9820
rect 67480 9818 67536 9820
rect 67240 9766 67286 9818
rect 67286 9766 67296 9818
rect 67320 9766 67350 9818
rect 67350 9766 67362 9818
rect 67362 9766 67376 9818
rect 67400 9766 67414 9818
rect 67414 9766 67426 9818
rect 67426 9766 67456 9818
rect 67480 9766 67490 9818
rect 67490 9766 67536 9818
rect 67240 9764 67296 9766
rect 67320 9764 67376 9766
rect 67400 9764 67456 9766
rect 67480 9764 67536 9766
rect 5140 9274 5196 9276
rect 5220 9274 5276 9276
rect 5300 9274 5356 9276
rect 5380 9274 5436 9276
rect 5140 9222 5186 9274
rect 5186 9222 5196 9274
rect 5220 9222 5250 9274
rect 5250 9222 5262 9274
rect 5262 9222 5276 9274
rect 5300 9222 5314 9274
rect 5314 9222 5326 9274
rect 5326 9222 5356 9274
rect 5380 9222 5390 9274
rect 5390 9222 5436 9274
rect 5140 9220 5196 9222
rect 5220 9220 5276 9222
rect 5300 9220 5356 9222
rect 5380 9220 5436 9222
rect 35860 9274 35916 9276
rect 35940 9274 35996 9276
rect 36020 9274 36076 9276
rect 36100 9274 36156 9276
rect 35860 9222 35906 9274
rect 35906 9222 35916 9274
rect 35940 9222 35970 9274
rect 35970 9222 35982 9274
rect 35982 9222 35996 9274
rect 36020 9222 36034 9274
rect 36034 9222 36046 9274
rect 36046 9222 36076 9274
rect 36100 9222 36110 9274
rect 36110 9222 36156 9274
rect 35860 9220 35916 9222
rect 35940 9220 35996 9222
rect 36020 9220 36076 9222
rect 36100 9220 36156 9222
rect 66580 9274 66636 9276
rect 66660 9274 66716 9276
rect 66740 9274 66796 9276
rect 66820 9274 66876 9276
rect 66580 9222 66626 9274
rect 66626 9222 66636 9274
rect 66660 9222 66690 9274
rect 66690 9222 66702 9274
rect 66702 9222 66716 9274
rect 66740 9222 66754 9274
rect 66754 9222 66766 9274
rect 66766 9222 66796 9274
rect 66820 9222 66830 9274
rect 66830 9222 66876 9274
rect 66580 9220 66636 9222
rect 66660 9220 66716 9222
rect 66740 9220 66796 9222
rect 66820 9220 66876 9222
rect 5800 8730 5856 8732
rect 5880 8730 5936 8732
rect 5960 8730 6016 8732
rect 6040 8730 6096 8732
rect 5800 8678 5846 8730
rect 5846 8678 5856 8730
rect 5880 8678 5910 8730
rect 5910 8678 5922 8730
rect 5922 8678 5936 8730
rect 5960 8678 5974 8730
rect 5974 8678 5986 8730
rect 5986 8678 6016 8730
rect 6040 8678 6050 8730
rect 6050 8678 6096 8730
rect 5800 8676 5856 8678
rect 5880 8676 5936 8678
rect 5960 8676 6016 8678
rect 6040 8676 6096 8678
rect 36520 8730 36576 8732
rect 36600 8730 36656 8732
rect 36680 8730 36736 8732
rect 36760 8730 36816 8732
rect 36520 8678 36566 8730
rect 36566 8678 36576 8730
rect 36600 8678 36630 8730
rect 36630 8678 36642 8730
rect 36642 8678 36656 8730
rect 36680 8678 36694 8730
rect 36694 8678 36706 8730
rect 36706 8678 36736 8730
rect 36760 8678 36770 8730
rect 36770 8678 36816 8730
rect 36520 8676 36576 8678
rect 36600 8676 36656 8678
rect 36680 8676 36736 8678
rect 36760 8676 36816 8678
rect 67240 8730 67296 8732
rect 67320 8730 67376 8732
rect 67400 8730 67456 8732
rect 67480 8730 67536 8732
rect 67240 8678 67286 8730
rect 67286 8678 67296 8730
rect 67320 8678 67350 8730
rect 67350 8678 67362 8730
rect 67362 8678 67376 8730
rect 67400 8678 67414 8730
rect 67414 8678 67426 8730
rect 67426 8678 67456 8730
rect 67480 8678 67490 8730
rect 67490 8678 67536 8730
rect 67240 8676 67296 8678
rect 67320 8676 67376 8678
rect 67400 8676 67456 8678
rect 67480 8676 67536 8678
rect 5140 8186 5196 8188
rect 5220 8186 5276 8188
rect 5300 8186 5356 8188
rect 5380 8186 5436 8188
rect 5140 8134 5186 8186
rect 5186 8134 5196 8186
rect 5220 8134 5250 8186
rect 5250 8134 5262 8186
rect 5262 8134 5276 8186
rect 5300 8134 5314 8186
rect 5314 8134 5326 8186
rect 5326 8134 5356 8186
rect 5380 8134 5390 8186
rect 5390 8134 5436 8186
rect 5140 8132 5196 8134
rect 5220 8132 5276 8134
rect 5300 8132 5356 8134
rect 5380 8132 5436 8134
rect 35860 8186 35916 8188
rect 35940 8186 35996 8188
rect 36020 8186 36076 8188
rect 36100 8186 36156 8188
rect 35860 8134 35906 8186
rect 35906 8134 35916 8186
rect 35940 8134 35970 8186
rect 35970 8134 35982 8186
rect 35982 8134 35996 8186
rect 36020 8134 36034 8186
rect 36034 8134 36046 8186
rect 36046 8134 36076 8186
rect 36100 8134 36110 8186
rect 36110 8134 36156 8186
rect 35860 8132 35916 8134
rect 35940 8132 35996 8134
rect 36020 8132 36076 8134
rect 36100 8132 36156 8134
rect 66580 8186 66636 8188
rect 66660 8186 66716 8188
rect 66740 8186 66796 8188
rect 66820 8186 66876 8188
rect 66580 8134 66626 8186
rect 66626 8134 66636 8186
rect 66660 8134 66690 8186
rect 66690 8134 66702 8186
rect 66702 8134 66716 8186
rect 66740 8134 66754 8186
rect 66754 8134 66766 8186
rect 66766 8134 66796 8186
rect 66820 8134 66830 8186
rect 66830 8134 66876 8186
rect 66580 8132 66636 8134
rect 66660 8132 66716 8134
rect 66740 8132 66796 8134
rect 66820 8132 66876 8134
rect 5800 7642 5856 7644
rect 5880 7642 5936 7644
rect 5960 7642 6016 7644
rect 6040 7642 6096 7644
rect 5800 7590 5846 7642
rect 5846 7590 5856 7642
rect 5880 7590 5910 7642
rect 5910 7590 5922 7642
rect 5922 7590 5936 7642
rect 5960 7590 5974 7642
rect 5974 7590 5986 7642
rect 5986 7590 6016 7642
rect 6040 7590 6050 7642
rect 6050 7590 6096 7642
rect 5800 7588 5856 7590
rect 5880 7588 5936 7590
rect 5960 7588 6016 7590
rect 6040 7588 6096 7590
rect 36520 7642 36576 7644
rect 36600 7642 36656 7644
rect 36680 7642 36736 7644
rect 36760 7642 36816 7644
rect 36520 7590 36566 7642
rect 36566 7590 36576 7642
rect 36600 7590 36630 7642
rect 36630 7590 36642 7642
rect 36642 7590 36656 7642
rect 36680 7590 36694 7642
rect 36694 7590 36706 7642
rect 36706 7590 36736 7642
rect 36760 7590 36770 7642
rect 36770 7590 36816 7642
rect 36520 7588 36576 7590
rect 36600 7588 36656 7590
rect 36680 7588 36736 7590
rect 36760 7588 36816 7590
rect 67240 7642 67296 7644
rect 67320 7642 67376 7644
rect 67400 7642 67456 7644
rect 67480 7642 67536 7644
rect 67240 7590 67286 7642
rect 67286 7590 67296 7642
rect 67320 7590 67350 7642
rect 67350 7590 67362 7642
rect 67362 7590 67376 7642
rect 67400 7590 67414 7642
rect 67414 7590 67426 7642
rect 67426 7590 67456 7642
rect 67480 7590 67490 7642
rect 67490 7590 67536 7642
rect 67240 7588 67296 7590
rect 67320 7588 67376 7590
rect 67400 7588 67456 7590
rect 67480 7588 67536 7590
rect 5140 7098 5196 7100
rect 5220 7098 5276 7100
rect 5300 7098 5356 7100
rect 5380 7098 5436 7100
rect 5140 7046 5186 7098
rect 5186 7046 5196 7098
rect 5220 7046 5250 7098
rect 5250 7046 5262 7098
rect 5262 7046 5276 7098
rect 5300 7046 5314 7098
rect 5314 7046 5326 7098
rect 5326 7046 5356 7098
rect 5380 7046 5390 7098
rect 5390 7046 5436 7098
rect 5140 7044 5196 7046
rect 5220 7044 5276 7046
rect 5300 7044 5356 7046
rect 5380 7044 5436 7046
rect 35860 7098 35916 7100
rect 35940 7098 35996 7100
rect 36020 7098 36076 7100
rect 36100 7098 36156 7100
rect 35860 7046 35906 7098
rect 35906 7046 35916 7098
rect 35940 7046 35970 7098
rect 35970 7046 35982 7098
rect 35982 7046 35996 7098
rect 36020 7046 36034 7098
rect 36034 7046 36046 7098
rect 36046 7046 36076 7098
rect 36100 7046 36110 7098
rect 36110 7046 36156 7098
rect 35860 7044 35916 7046
rect 35940 7044 35996 7046
rect 36020 7044 36076 7046
rect 36100 7044 36156 7046
rect 66580 7098 66636 7100
rect 66660 7098 66716 7100
rect 66740 7098 66796 7100
rect 66820 7098 66876 7100
rect 66580 7046 66626 7098
rect 66626 7046 66636 7098
rect 66660 7046 66690 7098
rect 66690 7046 66702 7098
rect 66702 7046 66716 7098
rect 66740 7046 66754 7098
rect 66754 7046 66766 7098
rect 66766 7046 66796 7098
rect 66820 7046 66830 7098
rect 66830 7046 66876 7098
rect 66580 7044 66636 7046
rect 66660 7044 66716 7046
rect 66740 7044 66796 7046
rect 66820 7044 66876 7046
rect 5800 6554 5856 6556
rect 5880 6554 5936 6556
rect 5960 6554 6016 6556
rect 6040 6554 6096 6556
rect 5800 6502 5846 6554
rect 5846 6502 5856 6554
rect 5880 6502 5910 6554
rect 5910 6502 5922 6554
rect 5922 6502 5936 6554
rect 5960 6502 5974 6554
rect 5974 6502 5986 6554
rect 5986 6502 6016 6554
rect 6040 6502 6050 6554
rect 6050 6502 6096 6554
rect 5800 6500 5856 6502
rect 5880 6500 5936 6502
rect 5960 6500 6016 6502
rect 6040 6500 6096 6502
rect 36520 6554 36576 6556
rect 36600 6554 36656 6556
rect 36680 6554 36736 6556
rect 36760 6554 36816 6556
rect 36520 6502 36566 6554
rect 36566 6502 36576 6554
rect 36600 6502 36630 6554
rect 36630 6502 36642 6554
rect 36642 6502 36656 6554
rect 36680 6502 36694 6554
rect 36694 6502 36706 6554
rect 36706 6502 36736 6554
rect 36760 6502 36770 6554
rect 36770 6502 36816 6554
rect 36520 6500 36576 6502
rect 36600 6500 36656 6502
rect 36680 6500 36736 6502
rect 36760 6500 36816 6502
rect 67240 6554 67296 6556
rect 67320 6554 67376 6556
rect 67400 6554 67456 6556
rect 67480 6554 67536 6556
rect 67240 6502 67286 6554
rect 67286 6502 67296 6554
rect 67320 6502 67350 6554
rect 67350 6502 67362 6554
rect 67362 6502 67376 6554
rect 67400 6502 67414 6554
rect 67414 6502 67426 6554
rect 67426 6502 67456 6554
rect 67480 6502 67490 6554
rect 67490 6502 67536 6554
rect 67240 6500 67296 6502
rect 67320 6500 67376 6502
rect 67400 6500 67456 6502
rect 67480 6500 67536 6502
rect 5140 6010 5196 6012
rect 5220 6010 5276 6012
rect 5300 6010 5356 6012
rect 5380 6010 5436 6012
rect 5140 5958 5186 6010
rect 5186 5958 5196 6010
rect 5220 5958 5250 6010
rect 5250 5958 5262 6010
rect 5262 5958 5276 6010
rect 5300 5958 5314 6010
rect 5314 5958 5326 6010
rect 5326 5958 5356 6010
rect 5380 5958 5390 6010
rect 5390 5958 5436 6010
rect 5140 5956 5196 5958
rect 5220 5956 5276 5958
rect 5300 5956 5356 5958
rect 5380 5956 5436 5958
rect 35860 6010 35916 6012
rect 35940 6010 35996 6012
rect 36020 6010 36076 6012
rect 36100 6010 36156 6012
rect 35860 5958 35906 6010
rect 35906 5958 35916 6010
rect 35940 5958 35970 6010
rect 35970 5958 35982 6010
rect 35982 5958 35996 6010
rect 36020 5958 36034 6010
rect 36034 5958 36046 6010
rect 36046 5958 36076 6010
rect 36100 5958 36110 6010
rect 36110 5958 36156 6010
rect 35860 5956 35916 5958
rect 35940 5956 35996 5958
rect 36020 5956 36076 5958
rect 36100 5956 36156 5958
rect 66580 6010 66636 6012
rect 66660 6010 66716 6012
rect 66740 6010 66796 6012
rect 66820 6010 66876 6012
rect 66580 5958 66626 6010
rect 66626 5958 66636 6010
rect 66660 5958 66690 6010
rect 66690 5958 66702 6010
rect 66702 5958 66716 6010
rect 66740 5958 66754 6010
rect 66754 5958 66766 6010
rect 66766 5958 66796 6010
rect 66820 5958 66830 6010
rect 66830 5958 66876 6010
rect 66580 5956 66636 5958
rect 66660 5956 66716 5958
rect 66740 5956 66796 5958
rect 66820 5956 66876 5958
rect 5800 5466 5856 5468
rect 5880 5466 5936 5468
rect 5960 5466 6016 5468
rect 6040 5466 6096 5468
rect 5800 5414 5846 5466
rect 5846 5414 5856 5466
rect 5880 5414 5910 5466
rect 5910 5414 5922 5466
rect 5922 5414 5936 5466
rect 5960 5414 5974 5466
rect 5974 5414 5986 5466
rect 5986 5414 6016 5466
rect 6040 5414 6050 5466
rect 6050 5414 6096 5466
rect 5800 5412 5856 5414
rect 5880 5412 5936 5414
rect 5960 5412 6016 5414
rect 6040 5412 6096 5414
rect 36520 5466 36576 5468
rect 36600 5466 36656 5468
rect 36680 5466 36736 5468
rect 36760 5466 36816 5468
rect 36520 5414 36566 5466
rect 36566 5414 36576 5466
rect 36600 5414 36630 5466
rect 36630 5414 36642 5466
rect 36642 5414 36656 5466
rect 36680 5414 36694 5466
rect 36694 5414 36706 5466
rect 36706 5414 36736 5466
rect 36760 5414 36770 5466
rect 36770 5414 36816 5466
rect 36520 5412 36576 5414
rect 36600 5412 36656 5414
rect 36680 5412 36736 5414
rect 36760 5412 36816 5414
rect 67240 5466 67296 5468
rect 67320 5466 67376 5468
rect 67400 5466 67456 5468
rect 67480 5466 67536 5468
rect 67240 5414 67286 5466
rect 67286 5414 67296 5466
rect 67320 5414 67350 5466
rect 67350 5414 67362 5466
rect 67362 5414 67376 5466
rect 67400 5414 67414 5466
rect 67414 5414 67426 5466
rect 67426 5414 67456 5466
rect 67480 5414 67490 5466
rect 67490 5414 67536 5466
rect 67240 5412 67296 5414
rect 67320 5412 67376 5414
rect 67400 5412 67456 5414
rect 67480 5412 67536 5414
rect 5140 4922 5196 4924
rect 5220 4922 5276 4924
rect 5300 4922 5356 4924
rect 5380 4922 5436 4924
rect 5140 4870 5186 4922
rect 5186 4870 5196 4922
rect 5220 4870 5250 4922
rect 5250 4870 5262 4922
rect 5262 4870 5276 4922
rect 5300 4870 5314 4922
rect 5314 4870 5326 4922
rect 5326 4870 5356 4922
rect 5380 4870 5390 4922
rect 5390 4870 5436 4922
rect 5140 4868 5196 4870
rect 5220 4868 5276 4870
rect 5300 4868 5356 4870
rect 5380 4868 5436 4870
rect 35860 4922 35916 4924
rect 35940 4922 35996 4924
rect 36020 4922 36076 4924
rect 36100 4922 36156 4924
rect 35860 4870 35906 4922
rect 35906 4870 35916 4922
rect 35940 4870 35970 4922
rect 35970 4870 35982 4922
rect 35982 4870 35996 4922
rect 36020 4870 36034 4922
rect 36034 4870 36046 4922
rect 36046 4870 36076 4922
rect 36100 4870 36110 4922
rect 36110 4870 36156 4922
rect 35860 4868 35916 4870
rect 35940 4868 35996 4870
rect 36020 4868 36076 4870
rect 36100 4868 36156 4870
rect 66580 4922 66636 4924
rect 66660 4922 66716 4924
rect 66740 4922 66796 4924
rect 66820 4922 66876 4924
rect 66580 4870 66626 4922
rect 66626 4870 66636 4922
rect 66660 4870 66690 4922
rect 66690 4870 66702 4922
rect 66702 4870 66716 4922
rect 66740 4870 66754 4922
rect 66754 4870 66766 4922
rect 66766 4870 66796 4922
rect 66820 4870 66830 4922
rect 66830 4870 66876 4922
rect 66580 4868 66636 4870
rect 66660 4868 66716 4870
rect 66740 4868 66796 4870
rect 66820 4868 66876 4870
rect 5800 4378 5856 4380
rect 5880 4378 5936 4380
rect 5960 4378 6016 4380
rect 6040 4378 6096 4380
rect 5800 4326 5846 4378
rect 5846 4326 5856 4378
rect 5880 4326 5910 4378
rect 5910 4326 5922 4378
rect 5922 4326 5936 4378
rect 5960 4326 5974 4378
rect 5974 4326 5986 4378
rect 5986 4326 6016 4378
rect 6040 4326 6050 4378
rect 6050 4326 6096 4378
rect 5800 4324 5856 4326
rect 5880 4324 5936 4326
rect 5960 4324 6016 4326
rect 6040 4324 6096 4326
rect 36520 4378 36576 4380
rect 36600 4378 36656 4380
rect 36680 4378 36736 4380
rect 36760 4378 36816 4380
rect 36520 4326 36566 4378
rect 36566 4326 36576 4378
rect 36600 4326 36630 4378
rect 36630 4326 36642 4378
rect 36642 4326 36656 4378
rect 36680 4326 36694 4378
rect 36694 4326 36706 4378
rect 36706 4326 36736 4378
rect 36760 4326 36770 4378
rect 36770 4326 36816 4378
rect 36520 4324 36576 4326
rect 36600 4324 36656 4326
rect 36680 4324 36736 4326
rect 36760 4324 36816 4326
rect 67240 4378 67296 4380
rect 67320 4378 67376 4380
rect 67400 4378 67456 4380
rect 67480 4378 67536 4380
rect 67240 4326 67286 4378
rect 67286 4326 67296 4378
rect 67320 4326 67350 4378
rect 67350 4326 67362 4378
rect 67362 4326 67376 4378
rect 67400 4326 67414 4378
rect 67414 4326 67426 4378
rect 67426 4326 67456 4378
rect 67480 4326 67490 4378
rect 67490 4326 67536 4378
rect 67240 4324 67296 4326
rect 67320 4324 67376 4326
rect 67400 4324 67456 4326
rect 67480 4324 67536 4326
rect 5140 3834 5196 3836
rect 5220 3834 5276 3836
rect 5300 3834 5356 3836
rect 5380 3834 5436 3836
rect 5140 3782 5186 3834
rect 5186 3782 5196 3834
rect 5220 3782 5250 3834
rect 5250 3782 5262 3834
rect 5262 3782 5276 3834
rect 5300 3782 5314 3834
rect 5314 3782 5326 3834
rect 5326 3782 5356 3834
rect 5380 3782 5390 3834
rect 5390 3782 5436 3834
rect 5140 3780 5196 3782
rect 5220 3780 5276 3782
rect 5300 3780 5356 3782
rect 5380 3780 5436 3782
rect 35860 3834 35916 3836
rect 35940 3834 35996 3836
rect 36020 3834 36076 3836
rect 36100 3834 36156 3836
rect 35860 3782 35906 3834
rect 35906 3782 35916 3834
rect 35940 3782 35970 3834
rect 35970 3782 35982 3834
rect 35982 3782 35996 3834
rect 36020 3782 36034 3834
rect 36034 3782 36046 3834
rect 36046 3782 36076 3834
rect 36100 3782 36110 3834
rect 36110 3782 36156 3834
rect 35860 3780 35916 3782
rect 35940 3780 35996 3782
rect 36020 3780 36076 3782
rect 36100 3780 36156 3782
rect 66580 3834 66636 3836
rect 66660 3834 66716 3836
rect 66740 3834 66796 3836
rect 66820 3834 66876 3836
rect 66580 3782 66626 3834
rect 66626 3782 66636 3834
rect 66660 3782 66690 3834
rect 66690 3782 66702 3834
rect 66702 3782 66716 3834
rect 66740 3782 66754 3834
rect 66754 3782 66766 3834
rect 66766 3782 66796 3834
rect 66820 3782 66830 3834
rect 66830 3782 66876 3834
rect 66580 3780 66636 3782
rect 66660 3780 66716 3782
rect 66740 3780 66796 3782
rect 66820 3780 66876 3782
rect 5800 3290 5856 3292
rect 5880 3290 5936 3292
rect 5960 3290 6016 3292
rect 6040 3290 6096 3292
rect 5800 3238 5846 3290
rect 5846 3238 5856 3290
rect 5880 3238 5910 3290
rect 5910 3238 5922 3290
rect 5922 3238 5936 3290
rect 5960 3238 5974 3290
rect 5974 3238 5986 3290
rect 5986 3238 6016 3290
rect 6040 3238 6050 3290
rect 6050 3238 6096 3290
rect 5800 3236 5856 3238
rect 5880 3236 5936 3238
rect 5960 3236 6016 3238
rect 6040 3236 6096 3238
rect 36520 3290 36576 3292
rect 36600 3290 36656 3292
rect 36680 3290 36736 3292
rect 36760 3290 36816 3292
rect 36520 3238 36566 3290
rect 36566 3238 36576 3290
rect 36600 3238 36630 3290
rect 36630 3238 36642 3290
rect 36642 3238 36656 3290
rect 36680 3238 36694 3290
rect 36694 3238 36706 3290
rect 36706 3238 36736 3290
rect 36760 3238 36770 3290
rect 36770 3238 36816 3290
rect 36520 3236 36576 3238
rect 36600 3236 36656 3238
rect 36680 3236 36736 3238
rect 36760 3236 36816 3238
rect 67240 3290 67296 3292
rect 67320 3290 67376 3292
rect 67400 3290 67456 3292
rect 67480 3290 67536 3292
rect 67240 3238 67286 3290
rect 67286 3238 67296 3290
rect 67320 3238 67350 3290
rect 67350 3238 67362 3290
rect 67362 3238 67376 3290
rect 67400 3238 67414 3290
rect 67414 3238 67426 3290
rect 67426 3238 67456 3290
rect 67480 3238 67490 3290
rect 67490 3238 67536 3290
rect 67240 3236 67296 3238
rect 67320 3236 67376 3238
rect 67400 3236 67456 3238
rect 67480 3236 67536 3238
rect 5140 2746 5196 2748
rect 5220 2746 5276 2748
rect 5300 2746 5356 2748
rect 5380 2746 5436 2748
rect 5140 2694 5186 2746
rect 5186 2694 5196 2746
rect 5220 2694 5250 2746
rect 5250 2694 5262 2746
rect 5262 2694 5276 2746
rect 5300 2694 5314 2746
rect 5314 2694 5326 2746
rect 5326 2694 5356 2746
rect 5380 2694 5390 2746
rect 5390 2694 5436 2746
rect 5140 2692 5196 2694
rect 5220 2692 5276 2694
rect 5300 2692 5356 2694
rect 5380 2692 5436 2694
rect 35860 2746 35916 2748
rect 35940 2746 35996 2748
rect 36020 2746 36076 2748
rect 36100 2746 36156 2748
rect 35860 2694 35906 2746
rect 35906 2694 35916 2746
rect 35940 2694 35970 2746
rect 35970 2694 35982 2746
rect 35982 2694 35996 2746
rect 36020 2694 36034 2746
rect 36034 2694 36046 2746
rect 36046 2694 36076 2746
rect 36100 2694 36110 2746
rect 36110 2694 36156 2746
rect 35860 2692 35916 2694
rect 35940 2692 35996 2694
rect 36020 2692 36076 2694
rect 36100 2692 36156 2694
rect 66580 2746 66636 2748
rect 66660 2746 66716 2748
rect 66740 2746 66796 2748
rect 66820 2746 66876 2748
rect 66580 2694 66626 2746
rect 66626 2694 66636 2746
rect 66660 2694 66690 2746
rect 66690 2694 66702 2746
rect 66702 2694 66716 2746
rect 66740 2694 66754 2746
rect 66754 2694 66766 2746
rect 66766 2694 66796 2746
rect 66820 2694 66830 2746
rect 66830 2694 66876 2746
rect 66580 2692 66636 2694
rect 66660 2692 66716 2694
rect 66740 2692 66796 2694
rect 66820 2692 66876 2694
rect 5800 2202 5856 2204
rect 5880 2202 5936 2204
rect 5960 2202 6016 2204
rect 6040 2202 6096 2204
rect 5800 2150 5846 2202
rect 5846 2150 5856 2202
rect 5880 2150 5910 2202
rect 5910 2150 5922 2202
rect 5922 2150 5936 2202
rect 5960 2150 5974 2202
rect 5974 2150 5986 2202
rect 5986 2150 6016 2202
rect 6040 2150 6050 2202
rect 6050 2150 6096 2202
rect 5800 2148 5856 2150
rect 5880 2148 5936 2150
rect 5960 2148 6016 2150
rect 6040 2148 6096 2150
rect 36520 2202 36576 2204
rect 36600 2202 36656 2204
rect 36680 2202 36736 2204
rect 36760 2202 36816 2204
rect 36520 2150 36566 2202
rect 36566 2150 36576 2202
rect 36600 2150 36630 2202
rect 36630 2150 36642 2202
rect 36642 2150 36656 2202
rect 36680 2150 36694 2202
rect 36694 2150 36706 2202
rect 36706 2150 36736 2202
rect 36760 2150 36770 2202
rect 36770 2150 36816 2202
rect 36520 2148 36576 2150
rect 36600 2148 36656 2150
rect 36680 2148 36736 2150
rect 36760 2148 36816 2150
rect 67240 2202 67296 2204
rect 67320 2202 67376 2204
rect 67400 2202 67456 2204
rect 67480 2202 67536 2204
rect 67240 2150 67286 2202
rect 67286 2150 67296 2202
rect 67320 2150 67350 2202
rect 67350 2150 67362 2202
rect 67362 2150 67376 2202
rect 67400 2150 67414 2202
rect 67414 2150 67426 2202
rect 67426 2150 67456 2202
rect 67480 2150 67490 2202
rect 67490 2150 67536 2202
rect 67240 2148 67296 2150
rect 67320 2148 67376 2150
rect 67400 2148 67456 2150
rect 67480 2148 67536 2150
<< metal3 >>
rect 5130 77824 5446 77825
rect 5130 77760 5136 77824
rect 5200 77760 5216 77824
rect 5280 77760 5296 77824
rect 5360 77760 5376 77824
rect 5440 77760 5446 77824
rect 5130 77759 5446 77760
rect 35850 77824 36166 77825
rect 35850 77760 35856 77824
rect 35920 77760 35936 77824
rect 36000 77760 36016 77824
rect 36080 77760 36096 77824
rect 36160 77760 36166 77824
rect 35850 77759 36166 77760
rect 66570 77824 66886 77825
rect 66570 77760 66576 77824
rect 66640 77760 66656 77824
rect 66720 77760 66736 77824
rect 66800 77760 66816 77824
rect 66880 77760 66886 77824
rect 66570 77759 66886 77760
rect 5790 77280 6106 77281
rect 5790 77216 5796 77280
rect 5860 77216 5876 77280
rect 5940 77216 5956 77280
rect 6020 77216 6036 77280
rect 6100 77216 6106 77280
rect 5790 77215 6106 77216
rect 36510 77280 36826 77281
rect 36510 77216 36516 77280
rect 36580 77216 36596 77280
rect 36660 77216 36676 77280
rect 36740 77216 36756 77280
rect 36820 77216 36826 77280
rect 36510 77215 36826 77216
rect 67230 77280 67546 77281
rect 67230 77216 67236 77280
rect 67300 77216 67316 77280
rect 67380 77216 67396 77280
rect 67460 77216 67476 77280
rect 67540 77216 67546 77280
rect 67230 77215 67546 77216
rect 5130 76736 5446 76737
rect 5130 76672 5136 76736
rect 5200 76672 5216 76736
rect 5280 76672 5296 76736
rect 5360 76672 5376 76736
rect 5440 76672 5446 76736
rect 5130 76671 5446 76672
rect 35850 76736 36166 76737
rect 35850 76672 35856 76736
rect 35920 76672 35936 76736
rect 36000 76672 36016 76736
rect 36080 76672 36096 76736
rect 36160 76672 36166 76736
rect 35850 76671 36166 76672
rect 66570 76736 66886 76737
rect 66570 76672 66576 76736
rect 66640 76672 66656 76736
rect 66720 76672 66736 76736
rect 66800 76672 66816 76736
rect 66880 76672 66886 76736
rect 66570 76671 66886 76672
rect 5790 76192 6106 76193
rect 5790 76128 5796 76192
rect 5860 76128 5876 76192
rect 5940 76128 5956 76192
rect 6020 76128 6036 76192
rect 6100 76128 6106 76192
rect 5790 76127 6106 76128
rect 36510 76192 36826 76193
rect 36510 76128 36516 76192
rect 36580 76128 36596 76192
rect 36660 76128 36676 76192
rect 36740 76128 36756 76192
rect 36820 76128 36826 76192
rect 36510 76127 36826 76128
rect 67230 76192 67546 76193
rect 67230 76128 67236 76192
rect 67300 76128 67316 76192
rect 67380 76128 67396 76192
rect 67460 76128 67476 76192
rect 67540 76128 67546 76192
rect 67230 76127 67546 76128
rect 5130 75648 5446 75649
rect 5130 75584 5136 75648
rect 5200 75584 5216 75648
rect 5280 75584 5296 75648
rect 5360 75584 5376 75648
rect 5440 75584 5446 75648
rect 5130 75583 5446 75584
rect 35850 75648 36166 75649
rect 35850 75584 35856 75648
rect 35920 75584 35936 75648
rect 36000 75584 36016 75648
rect 36080 75584 36096 75648
rect 36160 75584 36166 75648
rect 35850 75583 36166 75584
rect 66570 75648 66886 75649
rect 66570 75584 66576 75648
rect 66640 75584 66656 75648
rect 66720 75584 66736 75648
rect 66800 75584 66816 75648
rect 66880 75584 66886 75648
rect 66570 75583 66886 75584
rect 5790 75104 6106 75105
rect 5790 75040 5796 75104
rect 5860 75040 5876 75104
rect 5940 75040 5956 75104
rect 6020 75040 6036 75104
rect 6100 75040 6106 75104
rect 5790 75039 6106 75040
rect 36510 75104 36826 75105
rect 36510 75040 36516 75104
rect 36580 75040 36596 75104
rect 36660 75040 36676 75104
rect 36740 75040 36756 75104
rect 36820 75040 36826 75104
rect 36510 75039 36826 75040
rect 67230 75104 67546 75105
rect 67230 75040 67236 75104
rect 67300 75040 67316 75104
rect 67380 75040 67396 75104
rect 67460 75040 67476 75104
rect 67540 75040 67546 75104
rect 67230 75039 67546 75040
rect 5130 74560 5446 74561
rect 5130 74496 5136 74560
rect 5200 74496 5216 74560
rect 5280 74496 5296 74560
rect 5360 74496 5376 74560
rect 5440 74496 5446 74560
rect 5130 74495 5446 74496
rect 35850 74560 36166 74561
rect 35850 74496 35856 74560
rect 35920 74496 35936 74560
rect 36000 74496 36016 74560
rect 36080 74496 36096 74560
rect 36160 74496 36166 74560
rect 35850 74495 36166 74496
rect 66570 74560 66886 74561
rect 66570 74496 66576 74560
rect 66640 74496 66656 74560
rect 66720 74496 66736 74560
rect 66800 74496 66816 74560
rect 66880 74496 66886 74560
rect 66570 74495 66886 74496
rect 5790 74016 6106 74017
rect 5790 73952 5796 74016
rect 5860 73952 5876 74016
rect 5940 73952 5956 74016
rect 6020 73952 6036 74016
rect 6100 73952 6106 74016
rect 5790 73951 6106 73952
rect 36510 74016 36826 74017
rect 36510 73952 36516 74016
rect 36580 73952 36596 74016
rect 36660 73952 36676 74016
rect 36740 73952 36756 74016
rect 36820 73952 36826 74016
rect 36510 73951 36826 73952
rect 67230 74016 67546 74017
rect 67230 73952 67236 74016
rect 67300 73952 67316 74016
rect 67380 73952 67396 74016
rect 67460 73952 67476 74016
rect 67540 73952 67546 74016
rect 67230 73951 67546 73952
rect 5130 73472 5446 73473
rect 5130 73408 5136 73472
rect 5200 73408 5216 73472
rect 5280 73408 5296 73472
rect 5360 73408 5376 73472
rect 5440 73408 5446 73472
rect 5130 73407 5446 73408
rect 35850 73472 36166 73473
rect 35850 73408 35856 73472
rect 35920 73408 35936 73472
rect 36000 73408 36016 73472
rect 36080 73408 36096 73472
rect 36160 73408 36166 73472
rect 35850 73407 36166 73408
rect 66570 73472 66886 73473
rect 66570 73408 66576 73472
rect 66640 73408 66656 73472
rect 66720 73408 66736 73472
rect 66800 73408 66816 73472
rect 66880 73408 66886 73472
rect 66570 73407 66886 73408
rect 5790 72928 6106 72929
rect 5790 72864 5796 72928
rect 5860 72864 5876 72928
rect 5940 72864 5956 72928
rect 6020 72864 6036 72928
rect 6100 72864 6106 72928
rect 5790 72863 6106 72864
rect 36510 72928 36826 72929
rect 36510 72864 36516 72928
rect 36580 72864 36596 72928
rect 36660 72864 36676 72928
rect 36740 72864 36756 72928
rect 36820 72864 36826 72928
rect 36510 72863 36826 72864
rect 67230 72928 67546 72929
rect 67230 72864 67236 72928
rect 67300 72864 67316 72928
rect 67380 72864 67396 72928
rect 67460 72864 67476 72928
rect 67540 72864 67546 72928
rect 67230 72863 67546 72864
rect 5130 72384 5446 72385
rect 5130 72320 5136 72384
rect 5200 72320 5216 72384
rect 5280 72320 5296 72384
rect 5360 72320 5376 72384
rect 5440 72320 5446 72384
rect 5130 72319 5446 72320
rect 35850 72384 36166 72385
rect 35850 72320 35856 72384
rect 35920 72320 35936 72384
rect 36000 72320 36016 72384
rect 36080 72320 36096 72384
rect 36160 72320 36166 72384
rect 35850 72319 36166 72320
rect 66570 72384 66886 72385
rect 66570 72320 66576 72384
rect 66640 72320 66656 72384
rect 66720 72320 66736 72384
rect 66800 72320 66816 72384
rect 66880 72320 66886 72384
rect 66570 72319 66886 72320
rect 5790 71840 6106 71841
rect 5790 71776 5796 71840
rect 5860 71776 5876 71840
rect 5940 71776 5956 71840
rect 6020 71776 6036 71840
rect 6100 71776 6106 71840
rect 5790 71775 6106 71776
rect 36510 71840 36826 71841
rect 36510 71776 36516 71840
rect 36580 71776 36596 71840
rect 36660 71776 36676 71840
rect 36740 71776 36756 71840
rect 36820 71776 36826 71840
rect 36510 71775 36826 71776
rect 67230 71840 67546 71841
rect 67230 71776 67236 71840
rect 67300 71776 67316 71840
rect 67380 71776 67396 71840
rect 67460 71776 67476 71840
rect 67540 71776 67546 71840
rect 67230 71775 67546 71776
rect 5130 71296 5446 71297
rect 5130 71232 5136 71296
rect 5200 71232 5216 71296
rect 5280 71232 5296 71296
rect 5360 71232 5376 71296
rect 5440 71232 5446 71296
rect 5130 71231 5446 71232
rect 35850 71296 36166 71297
rect 35850 71232 35856 71296
rect 35920 71232 35936 71296
rect 36000 71232 36016 71296
rect 36080 71232 36096 71296
rect 36160 71232 36166 71296
rect 35850 71231 36166 71232
rect 66570 71296 66886 71297
rect 66570 71232 66576 71296
rect 66640 71232 66656 71296
rect 66720 71232 66736 71296
rect 66800 71232 66816 71296
rect 66880 71232 66886 71296
rect 66570 71231 66886 71232
rect 5790 70752 6106 70753
rect 5790 70688 5796 70752
rect 5860 70688 5876 70752
rect 5940 70688 5956 70752
rect 6020 70688 6036 70752
rect 6100 70688 6106 70752
rect 5790 70687 6106 70688
rect 36510 70752 36826 70753
rect 36510 70688 36516 70752
rect 36580 70688 36596 70752
rect 36660 70688 36676 70752
rect 36740 70688 36756 70752
rect 36820 70688 36826 70752
rect 36510 70687 36826 70688
rect 67230 70752 67546 70753
rect 67230 70688 67236 70752
rect 67300 70688 67316 70752
rect 67380 70688 67396 70752
rect 67460 70688 67476 70752
rect 67540 70688 67546 70752
rect 67230 70687 67546 70688
rect 5130 70208 5446 70209
rect 5130 70144 5136 70208
rect 5200 70144 5216 70208
rect 5280 70144 5296 70208
rect 5360 70144 5376 70208
rect 5440 70144 5446 70208
rect 5130 70143 5446 70144
rect 35850 70208 36166 70209
rect 35850 70144 35856 70208
rect 35920 70144 35936 70208
rect 36000 70144 36016 70208
rect 36080 70144 36096 70208
rect 36160 70144 36166 70208
rect 35850 70143 36166 70144
rect 66570 70208 66886 70209
rect 66570 70144 66576 70208
rect 66640 70144 66656 70208
rect 66720 70144 66736 70208
rect 66800 70144 66816 70208
rect 66880 70144 66886 70208
rect 66570 70143 66886 70144
rect 5790 69664 6106 69665
rect 5790 69600 5796 69664
rect 5860 69600 5876 69664
rect 5940 69600 5956 69664
rect 6020 69600 6036 69664
rect 6100 69600 6106 69664
rect 5790 69599 6106 69600
rect 36510 69664 36826 69665
rect 36510 69600 36516 69664
rect 36580 69600 36596 69664
rect 36660 69600 36676 69664
rect 36740 69600 36756 69664
rect 36820 69600 36826 69664
rect 36510 69599 36826 69600
rect 67230 69664 67546 69665
rect 67230 69600 67236 69664
rect 67300 69600 67316 69664
rect 67380 69600 67396 69664
rect 67460 69600 67476 69664
rect 67540 69600 67546 69664
rect 67230 69599 67546 69600
rect 5130 69120 5446 69121
rect 5130 69056 5136 69120
rect 5200 69056 5216 69120
rect 5280 69056 5296 69120
rect 5360 69056 5376 69120
rect 5440 69056 5446 69120
rect 5130 69055 5446 69056
rect 35850 69120 36166 69121
rect 35850 69056 35856 69120
rect 35920 69056 35936 69120
rect 36000 69056 36016 69120
rect 36080 69056 36096 69120
rect 36160 69056 36166 69120
rect 35850 69055 36166 69056
rect 66570 69120 66886 69121
rect 66570 69056 66576 69120
rect 66640 69056 66656 69120
rect 66720 69056 66736 69120
rect 66800 69056 66816 69120
rect 66880 69056 66886 69120
rect 66570 69055 66886 69056
rect 5790 68576 6106 68577
rect 5790 68512 5796 68576
rect 5860 68512 5876 68576
rect 5940 68512 5956 68576
rect 6020 68512 6036 68576
rect 6100 68512 6106 68576
rect 5790 68511 6106 68512
rect 36510 68576 36826 68577
rect 36510 68512 36516 68576
rect 36580 68512 36596 68576
rect 36660 68512 36676 68576
rect 36740 68512 36756 68576
rect 36820 68512 36826 68576
rect 36510 68511 36826 68512
rect 67230 68576 67546 68577
rect 67230 68512 67236 68576
rect 67300 68512 67316 68576
rect 67380 68512 67396 68576
rect 67460 68512 67476 68576
rect 67540 68512 67546 68576
rect 67230 68511 67546 68512
rect 5130 68032 5446 68033
rect 5130 67968 5136 68032
rect 5200 67968 5216 68032
rect 5280 67968 5296 68032
rect 5360 67968 5376 68032
rect 5440 67968 5446 68032
rect 5130 67967 5446 67968
rect 35850 68032 36166 68033
rect 35850 67968 35856 68032
rect 35920 67968 35936 68032
rect 36000 67968 36016 68032
rect 36080 67968 36096 68032
rect 36160 67968 36166 68032
rect 35850 67967 36166 67968
rect 66570 68032 66886 68033
rect 66570 67968 66576 68032
rect 66640 67968 66656 68032
rect 66720 67968 66736 68032
rect 66800 67968 66816 68032
rect 66880 67968 66886 68032
rect 66570 67967 66886 67968
rect 5790 67488 6106 67489
rect 5790 67424 5796 67488
rect 5860 67424 5876 67488
rect 5940 67424 5956 67488
rect 6020 67424 6036 67488
rect 6100 67424 6106 67488
rect 5790 67423 6106 67424
rect 36510 67488 36826 67489
rect 36510 67424 36516 67488
rect 36580 67424 36596 67488
rect 36660 67424 36676 67488
rect 36740 67424 36756 67488
rect 36820 67424 36826 67488
rect 36510 67423 36826 67424
rect 67230 67488 67546 67489
rect 67230 67424 67236 67488
rect 67300 67424 67316 67488
rect 67380 67424 67396 67488
rect 67460 67424 67476 67488
rect 67540 67424 67546 67488
rect 67230 67423 67546 67424
rect 5130 66944 5446 66945
rect 5130 66880 5136 66944
rect 5200 66880 5216 66944
rect 5280 66880 5296 66944
rect 5360 66880 5376 66944
rect 5440 66880 5446 66944
rect 5130 66879 5446 66880
rect 35850 66944 36166 66945
rect 35850 66880 35856 66944
rect 35920 66880 35936 66944
rect 36000 66880 36016 66944
rect 36080 66880 36096 66944
rect 36160 66880 36166 66944
rect 35850 66879 36166 66880
rect 66570 66944 66886 66945
rect 66570 66880 66576 66944
rect 66640 66880 66656 66944
rect 66720 66880 66736 66944
rect 66800 66880 66816 66944
rect 66880 66880 66886 66944
rect 66570 66879 66886 66880
rect 5790 66400 6106 66401
rect 5790 66336 5796 66400
rect 5860 66336 5876 66400
rect 5940 66336 5956 66400
rect 6020 66336 6036 66400
rect 6100 66336 6106 66400
rect 5790 66335 6106 66336
rect 36510 66400 36826 66401
rect 36510 66336 36516 66400
rect 36580 66336 36596 66400
rect 36660 66336 36676 66400
rect 36740 66336 36756 66400
rect 36820 66336 36826 66400
rect 36510 66335 36826 66336
rect 67230 66400 67546 66401
rect 67230 66336 67236 66400
rect 67300 66336 67316 66400
rect 67380 66336 67396 66400
rect 67460 66336 67476 66400
rect 67540 66336 67546 66400
rect 67230 66335 67546 66336
rect 5130 65856 5446 65857
rect 5130 65792 5136 65856
rect 5200 65792 5216 65856
rect 5280 65792 5296 65856
rect 5360 65792 5376 65856
rect 5440 65792 5446 65856
rect 5130 65791 5446 65792
rect 35850 65856 36166 65857
rect 35850 65792 35856 65856
rect 35920 65792 35936 65856
rect 36000 65792 36016 65856
rect 36080 65792 36096 65856
rect 36160 65792 36166 65856
rect 35850 65791 36166 65792
rect 66570 65856 66886 65857
rect 66570 65792 66576 65856
rect 66640 65792 66656 65856
rect 66720 65792 66736 65856
rect 66800 65792 66816 65856
rect 66880 65792 66886 65856
rect 66570 65791 66886 65792
rect 5790 65312 6106 65313
rect 5790 65248 5796 65312
rect 5860 65248 5876 65312
rect 5940 65248 5956 65312
rect 6020 65248 6036 65312
rect 6100 65248 6106 65312
rect 5790 65247 6106 65248
rect 36510 65312 36826 65313
rect 36510 65248 36516 65312
rect 36580 65248 36596 65312
rect 36660 65248 36676 65312
rect 36740 65248 36756 65312
rect 36820 65248 36826 65312
rect 36510 65247 36826 65248
rect 67230 65312 67546 65313
rect 67230 65248 67236 65312
rect 67300 65248 67316 65312
rect 67380 65248 67396 65312
rect 67460 65248 67476 65312
rect 67540 65248 67546 65312
rect 67230 65247 67546 65248
rect 5130 64768 5446 64769
rect 5130 64704 5136 64768
rect 5200 64704 5216 64768
rect 5280 64704 5296 64768
rect 5360 64704 5376 64768
rect 5440 64704 5446 64768
rect 5130 64703 5446 64704
rect 35850 64768 36166 64769
rect 35850 64704 35856 64768
rect 35920 64704 35936 64768
rect 36000 64704 36016 64768
rect 36080 64704 36096 64768
rect 36160 64704 36166 64768
rect 35850 64703 36166 64704
rect 66570 64768 66886 64769
rect 66570 64704 66576 64768
rect 66640 64704 66656 64768
rect 66720 64704 66736 64768
rect 66800 64704 66816 64768
rect 66880 64704 66886 64768
rect 66570 64703 66886 64704
rect 5790 64224 6106 64225
rect 5790 64160 5796 64224
rect 5860 64160 5876 64224
rect 5940 64160 5956 64224
rect 6020 64160 6036 64224
rect 6100 64160 6106 64224
rect 5790 64159 6106 64160
rect 36510 64224 36826 64225
rect 36510 64160 36516 64224
rect 36580 64160 36596 64224
rect 36660 64160 36676 64224
rect 36740 64160 36756 64224
rect 36820 64160 36826 64224
rect 36510 64159 36826 64160
rect 67230 64224 67546 64225
rect 67230 64160 67236 64224
rect 67300 64160 67316 64224
rect 67380 64160 67396 64224
rect 67460 64160 67476 64224
rect 67540 64160 67546 64224
rect 67230 64159 67546 64160
rect 5130 63680 5446 63681
rect 5130 63616 5136 63680
rect 5200 63616 5216 63680
rect 5280 63616 5296 63680
rect 5360 63616 5376 63680
rect 5440 63616 5446 63680
rect 5130 63615 5446 63616
rect 35850 63680 36166 63681
rect 35850 63616 35856 63680
rect 35920 63616 35936 63680
rect 36000 63616 36016 63680
rect 36080 63616 36096 63680
rect 36160 63616 36166 63680
rect 35850 63615 36166 63616
rect 66570 63680 66886 63681
rect 66570 63616 66576 63680
rect 66640 63616 66656 63680
rect 66720 63616 66736 63680
rect 66800 63616 66816 63680
rect 66880 63616 66886 63680
rect 66570 63615 66886 63616
rect 5790 63136 6106 63137
rect 5790 63072 5796 63136
rect 5860 63072 5876 63136
rect 5940 63072 5956 63136
rect 6020 63072 6036 63136
rect 6100 63072 6106 63136
rect 5790 63071 6106 63072
rect 36510 63136 36826 63137
rect 36510 63072 36516 63136
rect 36580 63072 36596 63136
rect 36660 63072 36676 63136
rect 36740 63072 36756 63136
rect 36820 63072 36826 63136
rect 36510 63071 36826 63072
rect 67230 63136 67546 63137
rect 67230 63072 67236 63136
rect 67300 63072 67316 63136
rect 67380 63072 67396 63136
rect 67460 63072 67476 63136
rect 67540 63072 67546 63136
rect 67230 63071 67546 63072
rect 5130 62592 5446 62593
rect 5130 62528 5136 62592
rect 5200 62528 5216 62592
rect 5280 62528 5296 62592
rect 5360 62528 5376 62592
rect 5440 62528 5446 62592
rect 5130 62527 5446 62528
rect 35850 62592 36166 62593
rect 35850 62528 35856 62592
rect 35920 62528 35936 62592
rect 36000 62528 36016 62592
rect 36080 62528 36096 62592
rect 36160 62528 36166 62592
rect 35850 62527 36166 62528
rect 66570 62592 66886 62593
rect 66570 62528 66576 62592
rect 66640 62528 66656 62592
rect 66720 62528 66736 62592
rect 66800 62528 66816 62592
rect 66880 62528 66886 62592
rect 66570 62527 66886 62528
rect 5790 62048 6106 62049
rect 5790 61984 5796 62048
rect 5860 61984 5876 62048
rect 5940 61984 5956 62048
rect 6020 61984 6036 62048
rect 6100 61984 6106 62048
rect 5790 61983 6106 61984
rect 36510 62048 36826 62049
rect 36510 61984 36516 62048
rect 36580 61984 36596 62048
rect 36660 61984 36676 62048
rect 36740 61984 36756 62048
rect 36820 61984 36826 62048
rect 36510 61983 36826 61984
rect 67230 62048 67546 62049
rect 67230 61984 67236 62048
rect 67300 61984 67316 62048
rect 67380 61984 67396 62048
rect 67460 61984 67476 62048
rect 67540 61984 67546 62048
rect 67230 61983 67546 61984
rect 5130 61504 5446 61505
rect 5130 61440 5136 61504
rect 5200 61440 5216 61504
rect 5280 61440 5296 61504
rect 5360 61440 5376 61504
rect 5440 61440 5446 61504
rect 5130 61439 5446 61440
rect 35850 61504 36166 61505
rect 35850 61440 35856 61504
rect 35920 61440 35936 61504
rect 36000 61440 36016 61504
rect 36080 61440 36096 61504
rect 36160 61440 36166 61504
rect 35850 61439 36166 61440
rect 66570 61504 66886 61505
rect 66570 61440 66576 61504
rect 66640 61440 66656 61504
rect 66720 61440 66736 61504
rect 66800 61440 66816 61504
rect 66880 61440 66886 61504
rect 66570 61439 66886 61440
rect 5790 60960 6106 60961
rect 5790 60896 5796 60960
rect 5860 60896 5876 60960
rect 5940 60896 5956 60960
rect 6020 60896 6036 60960
rect 6100 60896 6106 60960
rect 5790 60895 6106 60896
rect 36510 60960 36826 60961
rect 36510 60896 36516 60960
rect 36580 60896 36596 60960
rect 36660 60896 36676 60960
rect 36740 60896 36756 60960
rect 36820 60896 36826 60960
rect 36510 60895 36826 60896
rect 67230 60960 67546 60961
rect 67230 60896 67236 60960
rect 67300 60896 67316 60960
rect 67380 60896 67396 60960
rect 67460 60896 67476 60960
rect 67540 60896 67546 60960
rect 67230 60895 67546 60896
rect 5130 60416 5446 60417
rect 5130 60352 5136 60416
rect 5200 60352 5216 60416
rect 5280 60352 5296 60416
rect 5360 60352 5376 60416
rect 5440 60352 5446 60416
rect 5130 60351 5446 60352
rect 35850 60416 36166 60417
rect 35850 60352 35856 60416
rect 35920 60352 35936 60416
rect 36000 60352 36016 60416
rect 36080 60352 36096 60416
rect 36160 60352 36166 60416
rect 35850 60351 36166 60352
rect 66570 60416 66886 60417
rect 66570 60352 66576 60416
rect 66640 60352 66656 60416
rect 66720 60352 66736 60416
rect 66800 60352 66816 60416
rect 66880 60352 66886 60416
rect 66570 60351 66886 60352
rect 5790 59872 6106 59873
rect 5790 59808 5796 59872
rect 5860 59808 5876 59872
rect 5940 59808 5956 59872
rect 6020 59808 6036 59872
rect 6100 59808 6106 59872
rect 5790 59807 6106 59808
rect 36510 59872 36826 59873
rect 36510 59808 36516 59872
rect 36580 59808 36596 59872
rect 36660 59808 36676 59872
rect 36740 59808 36756 59872
rect 36820 59808 36826 59872
rect 36510 59807 36826 59808
rect 67230 59872 67546 59873
rect 67230 59808 67236 59872
rect 67300 59808 67316 59872
rect 67380 59808 67396 59872
rect 67460 59808 67476 59872
rect 67540 59808 67546 59872
rect 67230 59807 67546 59808
rect 5130 59328 5446 59329
rect 5130 59264 5136 59328
rect 5200 59264 5216 59328
rect 5280 59264 5296 59328
rect 5360 59264 5376 59328
rect 5440 59264 5446 59328
rect 5130 59263 5446 59264
rect 35850 59328 36166 59329
rect 35850 59264 35856 59328
rect 35920 59264 35936 59328
rect 36000 59264 36016 59328
rect 36080 59264 36096 59328
rect 36160 59264 36166 59328
rect 35850 59263 36166 59264
rect 66570 59328 66886 59329
rect 66570 59264 66576 59328
rect 66640 59264 66656 59328
rect 66720 59264 66736 59328
rect 66800 59264 66816 59328
rect 66880 59264 66886 59328
rect 66570 59263 66886 59264
rect 5790 58784 6106 58785
rect 5790 58720 5796 58784
rect 5860 58720 5876 58784
rect 5940 58720 5956 58784
rect 6020 58720 6036 58784
rect 6100 58720 6106 58784
rect 5790 58719 6106 58720
rect 36510 58784 36826 58785
rect 36510 58720 36516 58784
rect 36580 58720 36596 58784
rect 36660 58720 36676 58784
rect 36740 58720 36756 58784
rect 36820 58720 36826 58784
rect 36510 58719 36826 58720
rect 67230 58784 67546 58785
rect 67230 58720 67236 58784
rect 67300 58720 67316 58784
rect 67380 58720 67396 58784
rect 67460 58720 67476 58784
rect 67540 58720 67546 58784
rect 67230 58719 67546 58720
rect 5130 58240 5446 58241
rect 5130 58176 5136 58240
rect 5200 58176 5216 58240
rect 5280 58176 5296 58240
rect 5360 58176 5376 58240
rect 5440 58176 5446 58240
rect 5130 58175 5446 58176
rect 35850 58240 36166 58241
rect 35850 58176 35856 58240
rect 35920 58176 35936 58240
rect 36000 58176 36016 58240
rect 36080 58176 36096 58240
rect 36160 58176 36166 58240
rect 35850 58175 36166 58176
rect 66570 58240 66886 58241
rect 66570 58176 66576 58240
rect 66640 58176 66656 58240
rect 66720 58176 66736 58240
rect 66800 58176 66816 58240
rect 66880 58176 66886 58240
rect 66570 58175 66886 58176
rect 5790 57696 6106 57697
rect 5790 57632 5796 57696
rect 5860 57632 5876 57696
rect 5940 57632 5956 57696
rect 6020 57632 6036 57696
rect 6100 57632 6106 57696
rect 5790 57631 6106 57632
rect 36510 57696 36826 57697
rect 36510 57632 36516 57696
rect 36580 57632 36596 57696
rect 36660 57632 36676 57696
rect 36740 57632 36756 57696
rect 36820 57632 36826 57696
rect 36510 57631 36826 57632
rect 67230 57696 67546 57697
rect 67230 57632 67236 57696
rect 67300 57632 67316 57696
rect 67380 57632 67396 57696
rect 67460 57632 67476 57696
rect 67540 57632 67546 57696
rect 67230 57631 67546 57632
rect 5130 57152 5446 57153
rect 5130 57088 5136 57152
rect 5200 57088 5216 57152
rect 5280 57088 5296 57152
rect 5360 57088 5376 57152
rect 5440 57088 5446 57152
rect 5130 57087 5446 57088
rect 35850 57152 36166 57153
rect 35850 57088 35856 57152
rect 35920 57088 35936 57152
rect 36000 57088 36016 57152
rect 36080 57088 36096 57152
rect 36160 57088 36166 57152
rect 35850 57087 36166 57088
rect 66570 57152 66886 57153
rect 66570 57088 66576 57152
rect 66640 57088 66656 57152
rect 66720 57088 66736 57152
rect 66800 57088 66816 57152
rect 66880 57088 66886 57152
rect 66570 57087 66886 57088
rect 5790 56608 6106 56609
rect 5790 56544 5796 56608
rect 5860 56544 5876 56608
rect 5940 56544 5956 56608
rect 6020 56544 6036 56608
rect 6100 56544 6106 56608
rect 5790 56543 6106 56544
rect 36510 56608 36826 56609
rect 36510 56544 36516 56608
rect 36580 56544 36596 56608
rect 36660 56544 36676 56608
rect 36740 56544 36756 56608
rect 36820 56544 36826 56608
rect 36510 56543 36826 56544
rect 67230 56608 67546 56609
rect 67230 56544 67236 56608
rect 67300 56544 67316 56608
rect 67380 56544 67396 56608
rect 67460 56544 67476 56608
rect 67540 56544 67546 56608
rect 67230 56543 67546 56544
rect 5130 56064 5446 56065
rect 5130 56000 5136 56064
rect 5200 56000 5216 56064
rect 5280 56000 5296 56064
rect 5360 56000 5376 56064
rect 5440 56000 5446 56064
rect 5130 55999 5446 56000
rect 35850 56064 36166 56065
rect 35850 56000 35856 56064
rect 35920 56000 35936 56064
rect 36000 56000 36016 56064
rect 36080 56000 36096 56064
rect 36160 56000 36166 56064
rect 35850 55999 36166 56000
rect 66570 56064 66886 56065
rect 66570 56000 66576 56064
rect 66640 56000 66656 56064
rect 66720 56000 66736 56064
rect 66800 56000 66816 56064
rect 66880 56000 66886 56064
rect 66570 55999 66886 56000
rect 5790 55520 6106 55521
rect 5790 55456 5796 55520
rect 5860 55456 5876 55520
rect 5940 55456 5956 55520
rect 6020 55456 6036 55520
rect 6100 55456 6106 55520
rect 5790 55455 6106 55456
rect 36510 55520 36826 55521
rect 36510 55456 36516 55520
rect 36580 55456 36596 55520
rect 36660 55456 36676 55520
rect 36740 55456 36756 55520
rect 36820 55456 36826 55520
rect 36510 55455 36826 55456
rect 67230 55520 67546 55521
rect 67230 55456 67236 55520
rect 67300 55456 67316 55520
rect 67380 55456 67396 55520
rect 67460 55456 67476 55520
rect 67540 55456 67546 55520
rect 67230 55455 67546 55456
rect 5130 54976 5446 54977
rect 5130 54912 5136 54976
rect 5200 54912 5216 54976
rect 5280 54912 5296 54976
rect 5360 54912 5376 54976
rect 5440 54912 5446 54976
rect 5130 54911 5446 54912
rect 35850 54976 36166 54977
rect 35850 54912 35856 54976
rect 35920 54912 35936 54976
rect 36000 54912 36016 54976
rect 36080 54912 36096 54976
rect 36160 54912 36166 54976
rect 35850 54911 36166 54912
rect 66570 54976 66886 54977
rect 66570 54912 66576 54976
rect 66640 54912 66656 54976
rect 66720 54912 66736 54976
rect 66800 54912 66816 54976
rect 66880 54912 66886 54976
rect 66570 54911 66886 54912
rect 5790 54432 6106 54433
rect 5790 54368 5796 54432
rect 5860 54368 5876 54432
rect 5940 54368 5956 54432
rect 6020 54368 6036 54432
rect 6100 54368 6106 54432
rect 5790 54367 6106 54368
rect 36510 54432 36826 54433
rect 36510 54368 36516 54432
rect 36580 54368 36596 54432
rect 36660 54368 36676 54432
rect 36740 54368 36756 54432
rect 36820 54368 36826 54432
rect 36510 54367 36826 54368
rect 67230 54432 67546 54433
rect 67230 54368 67236 54432
rect 67300 54368 67316 54432
rect 67380 54368 67396 54432
rect 67460 54368 67476 54432
rect 67540 54368 67546 54432
rect 67230 54367 67546 54368
rect 5130 53888 5446 53889
rect 5130 53824 5136 53888
rect 5200 53824 5216 53888
rect 5280 53824 5296 53888
rect 5360 53824 5376 53888
rect 5440 53824 5446 53888
rect 5130 53823 5446 53824
rect 35850 53888 36166 53889
rect 35850 53824 35856 53888
rect 35920 53824 35936 53888
rect 36000 53824 36016 53888
rect 36080 53824 36096 53888
rect 36160 53824 36166 53888
rect 35850 53823 36166 53824
rect 66570 53888 66886 53889
rect 66570 53824 66576 53888
rect 66640 53824 66656 53888
rect 66720 53824 66736 53888
rect 66800 53824 66816 53888
rect 66880 53824 66886 53888
rect 66570 53823 66886 53824
rect 5790 53344 6106 53345
rect 5790 53280 5796 53344
rect 5860 53280 5876 53344
rect 5940 53280 5956 53344
rect 6020 53280 6036 53344
rect 6100 53280 6106 53344
rect 5790 53279 6106 53280
rect 36510 53344 36826 53345
rect 36510 53280 36516 53344
rect 36580 53280 36596 53344
rect 36660 53280 36676 53344
rect 36740 53280 36756 53344
rect 36820 53280 36826 53344
rect 36510 53279 36826 53280
rect 67230 53344 67546 53345
rect 67230 53280 67236 53344
rect 67300 53280 67316 53344
rect 67380 53280 67396 53344
rect 67460 53280 67476 53344
rect 67540 53280 67546 53344
rect 67230 53279 67546 53280
rect 5130 52800 5446 52801
rect 5130 52736 5136 52800
rect 5200 52736 5216 52800
rect 5280 52736 5296 52800
rect 5360 52736 5376 52800
rect 5440 52736 5446 52800
rect 5130 52735 5446 52736
rect 35850 52800 36166 52801
rect 35850 52736 35856 52800
rect 35920 52736 35936 52800
rect 36000 52736 36016 52800
rect 36080 52736 36096 52800
rect 36160 52736 36166 52800
rect 35850 52735 36166 52736
rect 66570 52800 66886 52801
rect 66570 52736 66576 52800
rect 66640 52736 66656 52800
rect 66720 52736 66736 52800
rect 66800 52736 66816 52800
rect 66880 52736 66886 52800
rect 66570 52735 66886 52736
rect 5790 52256 6106 52257
rect 5790 52192 5796 52256
rect 5860 52192 5876 52256
rect 5940 52192 5956 52256
rect 6020 52192 6036 52256
rect 6100 52192 6106 52256
rect 5790 52191 6106 52192
rect 36510 52256 36826 52257
rect 36510 52192 36516 52256
rect 36580 52192 36596 52256
rect 36660 52192 36676 52256
rect 36740 52192 36756 52256
rect 36820 52192 36826 52256
rect 36510 52191 36826 52192
rect 67230 52256 67546 52257
rect 67230 52192 67236 52256
rect 67300 52192 67316 52256
rect 67380 52192 67396 52256
rect 67460 52192 67476 52256
rect 67540 52192 67546 52256
rect 67230 52191 67546 52192
rect 77569 51778 77635 51781
rect 79200 51778 80000 51808
rect 77569 51776 80000 51778
rect 77569 51720 77574 51776
rect 77630 51720 80000 51776
rect 77569 51718 80000 51720
rect 77569 51715 77635 51718
rect 5130 51712 5446 51713
rect 5130 51648 5136 51712
rect 5200 51648 5216 51712
rect 5280 51648 5296 51712
rect 5360 51648 5376 51712
rect 5440 51648 5446 51712
rect 5130 51647 5446 51648
rect 35850 51712 36166 51713
rect 35850 51648 35856 51712
rect 35920 51648 35936 51712
rect 36000 51648 36016 51712
rect 36080 51648 36096 51712
rect 36160 51648 36166 51712
rect 35850 51647 36166 51648
rect 66570 51712 66886 51713
rect 66570 51648 66576 51712
rect 66640 51648 66656 51712
rect 66720 51648 66736 51712
rect 66800 51648 66816 51712
rect 66880 51648 66886 51712
rect 79200 51688 80000 51718
rect 66570 51647 66886 51648
rect 5790 51168 6106 51169
rect 5790 51104 5796 51168
rect 5860 51104 5876 51168
rect 5940 51104 5956 51168
rect 6020 51104 6036 51168
rect 6100 51104 6106 51168
rect 5790 51103 6106 51104
rect 36510 51168 36826 51169
rect 36510 51104 36516 51168
rect 36580 51104 36596 51168
rect 36660 51104 36676 51168
rect 36740 51104 36756 51168
rect 36820 51104 36826 51168
rect 36510 51103 36826 51104
rect 67230 51168 67546 51169
rect 67230 51104 67236 51168
rect 67300 51104 67316 51168
rect 67380 51104 67396 51168
rect 67460 51104 67476 51168
rect 67540 51104 67546 51168
rect 67230 51103 67546 51104
rect 5130 50624 5446 50625
rect 5130 50560 5136 50624
rect 5200 50560 5216 50624
rect 5280 50560 5296 50624
rect 5360 50560 5376 50624
rect 5440 50560 5446 50624
rect 5130 50559 5446 50560
rect 35850 50624 36166 50625
rect 35850 50560 35856 50624
rect 35920 50560 35936 50624
rect 36000 50560 36016 50624
rect 36080 50560 36096 50624
rect 36160 50560 36166 50624
rect 35850 50559 36166 50560
rect 66570 50624 66886 50625
rect 66570 50560 66576 50624
rect 66640 50560 66656 50624
rect 66720 50560 66736 50624
rect 66800 50560 66816 50624
rect 66880 50560 66886 50624
rect 66570 50559 66886 50560
rect 5790 50080 6106 50081
rect 5790 50016 5796 50080
rect 5860 50016 5876 50080
rect 5940 50016 5956 50080
rect 6020 50016 6036 50080
rect 6100 50016 6106 50080
rect 5790 50015 6106 50016
rect 36510 50080 36826 50081
rect 36510 50016 36516 50080
rect 36580 50016 36596 50080
rect 36660 50016 36676 50080
rect 36740 50016 36756 50080
rect 36820 50016 36826 50080
rect 36510 50015 36826 50016
rect 67230 50080 67546 50081
rect 67230 50016 67236 50080
rect 67300 50016 67316 50080
rect 67380 50016 67396 50080
rect 67460 50016 67476 50080
rect 67540 50016 67546 50080
rect 67230 50015 67546 50016
rect 77569 49738 77635 49741
rect 79200 49738 80000 49768
rect 77569 49736 80000 49738
rect 77569 49680 77574 49736
rect 77630 49680 80000 49736
rect 77569 49678 80000 49680
rect 77569 49675 77635 49678
rect 79200 49648 80000 49678
rect 5130 49536 5446 49537
rect 5130 49472 5136 49536
rect 5200 49472 5216 49536
rect 5280 49472 5296 49536
rect 5360 49472 5376 49536
rect 5440 49472 5446 49536
rect 5130 49471 5446 49472
rect 35850 49536 36166 49537
rect 35850 49472 35856 49536
rect 35920 49472 35936 49536
rect 36000 49472 36016 49536
rect 36080 49472 36096 49536
rect 36160 49472 36166 49536
rect 35850 49471 36166 49472
rect 66570 49536 66886 49537
rect 66570 49472 66576 49536
rect 66640 49472 66656 49536
rect 66720 49472 66736 49536
rect 66800 49472 66816 49536
rect 66880 49472 66886 49536
rect 66570 49471 66886 49472
rect 5790 48992 6106 48993
rect 5790 48928 5796 48992
rect 5860 48928 5876 48992
rect 5940 48928 5956 48992
rect 6020 48928 6036 48992
rect 6100 48928 6106 48992
rect 5790 48927 6106 48928
rect 36510 48992 36826 48993
rect 36510 48928 36516 48992
rect 36580 48928 36596 48992
rect 36660 48928 36676 48992
rect 36740 48928 36756 48992
rect 36820 48928 36826 48992
rect 36510 48927 36826 48928
rect 67230 48992 67546 48993
rect 67230 48928 67236 48992
rect 67300 48928 67316 48992
rect 67380 48928 67396 48992
rect 67460 48928 67476 48992
rect 67540 48928 67546 48992
rect 67230 48927 67546 48928
rect 5130 48448 5446 48449
rect 5130 48384 5136 48448
rect 5200 48384 5216 48448
rect 5280 48384 5296 48448
rect 5360 48384 5376 48448
rect 5440 48384 5446 48448
rect 5130 48383 5446 48384
rect 35850 48448 36166 48449
rect 35850 48384 35856 48448
rect 35920 48384 35936 48448
rect 36000 48384 36016 48448
rect 36080 48384 36096 48448
rect 36160 48384 36166 48448
rect 35850 48383 36166 48384
rect 66570 48448 66886 48449
rect 66570 48384 66576 48448
rect 66640 48384 66656 48448
rect 66720 48384 66736 48448
rect 66800 48384 66816 48448
rect 66880 48384 66886 48448
rect 66570 48383 66886 48384
rect 5790 47904 6106 47905
rect 5790 47840 5796 47904
rect 5860 47840 5876 47904
rect 5940 47840 5956 47904
rect 6020 47840 6036 47904
rect 6100 47840 6106 47904
rect 5790 47839 6106 47840
rect 36510 47904 36826 47905
rect 36510 47840 36516 47904
rect 36580 47840 36596 47904
rect 36660 47840 36676 47904
rect 36740 47840 36756 47904
rect 36820 47840 36826 47904
rect 36510 47839 36826 47840
rect 67230 47904 67546 47905
rect 67230 47840 67236 47904
rect 67300 47840 67316 47904
rect 67380 47840 67396 47904
rect 67460 47840 67476 47904
rect 67540 47840 67546 47904
rect 67230 47839 67546 47840
rect 5130 47360 5446 47361
rect 5130 47296 5136 47360
rect 5200 47296 5216 47360
rect 5280 47296 5296 47360
rect 5360 47296 5376 47360
rect 5440 47296 5446 47360
rect 5130 47295 5446 47296
rect 35850 47360 36166 47361
rect 35850 47296 35856 47360
rect 35920 47296 35936 47360
rect 36000 47296 36016 47360
rect 36080 47296 36096 47360
rect 36160 47296 36166 47360
rect 35850 47295 36166 47296
rect 66570 47360 66886 47361
rect 66570 47296 66576 47360
rect 66640 47296 66656 47360
rect 66720 47296 66736 47360
rect 66800 47296 66816 47360
rect 66880 47296 66886 47360
rect 66570 47295 66886 47296
rect 5790 46816 6106 46817
rect 5790 46752 5796 46816
rect 5860 46752 5876 46816
rect 5940 46752 5956 46816
rect 6020 46752 6036 46816
rect 6100 46752 6106 46816
rect 5790 46751 6106 46752
rect 36510 46816 36826 46817
rect 36510 46752 36516 46816
rect 36580 46752 36596 46816
rect 36660 46752 36676 46816
rect 36740 46752 36756 46816
rect 36820 46752 36826 46816
rect 36510 46751 36826 46752
rect 67230 46816 67546 46817
rect 67230 46752 67236 46816
rect 67300 46752 67316 46816
rect 67380 46752 67396 46816
rect 67460 46752 67476 46816
rect 67540 46752 67546 46816
rect 67230 46751 67546 46752
rect 5130 46272 5446 46273
rect 5130 46208 5136 46272
rect 5200 46208 5216 46272
rect 5280 46208 5296 46272
rect 5360 46208 5376 46272
rect 5440 46208 5446 46272
rect 5130 46207 5446 46208
rect 35850 46272 36166 46273
rect 35850 46208 35856 46272
rect 35920 46208 35936 46272
rect 36000 46208 36016 46272
rect 36080 46208 36096 46272
rect 36160 46208 36166 46272
rect 35850 46207 36166 46208
rect 66570 46272 66886 46273
rect 66570 46208 66576 46272
rect 66640 46208 66656 46272
rect 66720 46208 66736 46272
rect 66800 46208 66816 46272
rect 66880 46208 66886 46272
rect 66570 46207 66886 46208
rect 5790 45728 6106 45729
rect 0 45658 800 45688
rect 5790 45664 5796 45728
rect 5860 45664 5876 45728
rect 5940 45664 5956 45728
rect 6020 45664 6036 45728
rect 6100 45664 6106 45728
rect 5790 45663 6106 45664
rect 36510 45728 36826 45729
rect 36510 45664 36516 45728
rect 36580 45664 36596 45728
rect 36660 45664 36676 45728
rect 36740 45664 36756 45728
rect 36820 45664 36826 45728
rect 36510 45663 36826 45664
rect 67230 45728 67546 45729
rect 67230 45664 67236 45728
rect 67300 45664 67316 45728
rect 67380 45664 67396 45728
rect 67460 45664 67476 45728
rect 67540 45664 67546 45728
rect 67230 45663 67546 45664
rect 1301 45658 1367 45661
rect 0 45656 1367 45658
rect 0 45600 1306 45656
rect 1362 45600 1367 45656
rect 0 45598 1367 45600
rect 0 45568 800 45598
rect 1301 45595 1367 45598
rect 5130 45184 5446 45185
rect 5130 45120 5136 45184
rect 5200 45120 5216 45184
rect 5280 45120 5296 45184
rect 5360 45120 5376 45184
rect 5440 45120 5446 45184
rect 5130 45119 5446 45120
rect 35850 45184 36166 45185
rect 35850 45120 35856 45184
rect 35920 45120 35936 45184
rect 36000 45120 36016 45184
rect 36080 45120 36096 45184
rect 36160 45120 36166 45184
rect 35850 45119 36166 45120
rect 66570 45184 66886 45185
rect 66570 45120 66576 45184
rect 66640 45120 66656 45184
rect 66720 45120 66736 45184
rect 66800 45120 66816 45184
rect 66880 45120 66886 45184
rect 66570 45119 66886 45120
rect 5790 44640 6106 44641
rect 5790 44576 5796 44640
rect 5860 44576 5876 44640
rect 5940 44576 5956 44640
rect 6020 44576 6036 44640
rect 6100 44576 6106 44640
rect 5790 44575 6106 44576
rect 36510 44640 36826 44641
rect 36510 44576 36516 44640
rect 36580 44576 36596 44640
rect 36660 44576 36676 44640
rect 36740 44576 36756 44640
rect 36820 44576 36826 44640
rect 36510 44575 36826 44576
rect 67230 44640 67546 44641
rect 67230 44576 67236 44640
rect 67300 44576 67316 44640
rect 67380 44576 67396 44640
rect 67460 44576 67476 44640
rect 67540 44576 67546 44640
rect 67230 44575 67546 44576
rect 5130 44096 5446 44097
rect 5130 44032 5136 44096
rect 5200 44032 5216 44096
rect 5280 44032 5296 44096
rect 5360 44032 5376 44096
rect 5440 44032 5446 44096
rect 5130 44031 5446 44032
rect 35850 44096 36166 44097
rect 35850 44032 35856 44096
rect 35920 44032 35936 44096
rect 36000 44032 36016 44096
rect 36080 44032 36096 44096
rect 36160 44032 36166 44096
rect 35850 44031 36166 44032
rect 66570 44096 66886 44097
rect 66570 44032 66576 44096
rect 66640 44032 66656 44096
rect 66720 44032 66736 44096
rect 66800 44032 66816 44096
rect 66880 44032 66886 44096
rect 66570 44031 66886 44032
rect 5790 43552 6106 43553
rect 5790 43488 5796 43552
rect 5860 43488 5876 43552
rect 5940 43488 5956 43552
rect 6020 43488 6036 43552
rect 6100 43488 6106 43552
rect 5790 43487 6106 43488
rect 36510 43552 36826 43553
rect 36510 43488 36516 43552
rect 36580 43488 36596 43552
rect 36660 43488 36676 43552
rect 36740 43488 36756 43552
rect 36820 43488 36826 43552
rect 36510 43487 36826 43488
rect 67230 43552 67546 43553
rect 67230 43488 67236 43552
rect 67300 43488 67316 43552
rect 67380 43488 67396 43552
rect 67460 43488 67476 43552
rect 67540 43488 67546 43552
rect 67230 43487 67546 43488
rect 5130 43008 5446 43009
rect 5130 42944 5136 43008
rect 5200 42944 5216 43008
rect 5280 42944 5296 43008
rect 5360 42944 5376 43008
rect 5440 42944 5446 43008
rect 5130 42943 5446 42944
rect 35850 43008 36166 43009
rect 35850 42944 35856 43008
rect 35920 42944 35936 43008
rect 36000 42944 36016 43008
rect 36080 42944 36096 43008
rect 36160 42944 36166 43008
rect 35850 42943 36166 42944
rect 66570 43008 66886 43009
rect 66570 42944 66576 43008
rect 66640 42944 66656 43008
rect 66720 42944 66736 43008
rect 66800 42944 66816 43008
rect 66880 42944 66886 43008
rect 66570 42943 66886 42944
rect 5790 42464 6106 42465
rect 5790 42400 5796 42464
rect 5860 42400 5876 42464
rect 5940 42400 5956 42464
rect 6020 42400 6036 42464
rect 6100 42400 6106 42464
rect 5790 42399 6106 42400
rect 36510 42464 36826 42465
rect 36510 42400 36516 42464
rect 36580 42400 36596 42464
rect 36660 42400 36676 42464
rect 36740 42400 36756 42464
rect 36820 42400 36826 42464
rect 36510 42399 36826 42400
rect 67230 42464 67546 42465
rect 67230 42400 67236 42464
rect 67300 42400 67316 42464
rect 67380 42400 67396 42464
rect 67460 42400 67476 42464
rect 67540 42400 67546 42464
rect 67230 42399 67546 42400
rect 5130 41920 5446 41921
rect 5130 41856 5136 41920
rect 5200 41856 5216 41920
rect 5280 41856 5296 41920
rect 5360 41856 5376 41920
rect 5440 41856 5446 41920
rect 5130 41855 5446 41856
rect 35850 41920 36166 41921
rect 35850 41856 35856 41920
rect 35920 41856 35936 41920
rect 36000 41856 36016 41920
rect 36080 41856 36096 41920
rect 36160 41856 36166 41920
rect 35850 41855 36166 41856
rect 66570 41920 66886 41921
rect 66570 41856 66576 41920
rect 66640 41856 66656 41920
rect 66720 41856 66736 41920
rect 66800 41856 66816 41920
rect 66880 41856 66886 41920
rect 66570 41855 66886 41856
rect 0 41578 800 41608
rect 1209 41578 1275 41581
rect 0 41576 1275 41578
rect 0 41520 1214 41576
rect 1270 41520 1275 41576
rect 0 41518 1275 41520
rect 0 41488 800 41518
rect 1209 41515 1275 41518
rect 5790 41376 6106 41377
rect 5790 41312 5796 41376
rect 5860 41312 5876 41376
rect 5940 41312 5956 41376
rect 6020 41312 6036 41376
rect 6100 41312 6106 41376
rect 5790 41311 6106 41312
rect 36510 41376 36826 41377
rect 36510 41312 36516 41376
rect 36580 41312 36596 41376
rect 36660 41312 36676 41376
rect 36740 41312 36756 41376
rect 36820 41312 36826 41376
rect 36510 41311 36826 41312
rect 67230 41376 67546 41377
rect 67230 41312 67236 41376
rect 67300 41312 67316 41376
rect 67380 41312 67396 41376
rect 67460 41312 67476 41376
rect 67540 41312 67546 41376
rect 67230 41311 67546 41312
rect 5130 40832 5446 40833
rect 5130 40768 5136 40832
rect 5200 40768 5216 40832
rect 5280 40768 5296 40832
rect 5360 40768 5376 40832
rect 5440 40768 5446 40832
rect 5130 40767 5446 40768
rect 35850 40832 36166 40833
rect 35850 40768 35856 40832
rect 35920 40768 35936 40832
rect 36000 40768 36016 40832
rect 36080 40768 36096 40832
rect 36160 40768 36166 40832
rect 35850 40767 36166 40768
rect 66570 40832 66886 40833
rect 66570 40768 66576 40832
rect 66640 40768 66656 40832
rect 66720 40768 66736 40832
rect 66800 40768 66816 40832
rect 66880 40768 66886 40832
rect 66570 40767 66886 40768
rect 5790 40288 6106 40289
rect 5790 40224 5796 40288
rect 5860 40224 5876 40288
rect 5940 40224 5956 40288
rect 6020 40224 6036 40288
rect 6100 40224 6106 40288
rect 5790 40223 6106 40224
rect 36510 40288 36826 40289
rect 36510 40224 36516 40288
rect 36580 40224 36596 40288
rect 36660 40224 36676 40288
rect 36740 40224 36756 40288
rect 36820 40224 36826 40288
rect 36510 40223 36826 40224
rect 67230 40288 67546 40289
rect 67230 40224 67236 40288
rect 67300 40224 67316 40288
rect 67380 40224 67396 40288
rect 67460 40224 67476 40288
rect 67540 40224 67546 40288
rect 67230 40223 67546 40224
rect 5130 39744 5446 39745
rect 5130 39680 5136 39744
rect 5200 39680 5216 39744
rect 5280 39680 5296 39744
rect 5360 39680 5376 39744
rect 5440 39680 5446 39744
rect 5130 39679 5446 39680
rect 35850 39744 36166 39745
rect 35850 39680 35856 39744
rect 35920 39680 35936 39744
rect 36000 39680 36016 39744
rect 36080 39680 36096 39744
rect 36160 39680 36166 39744
rect 35850 39679 36166 39680
rect 66570 39744 66886 39745
rect 66570 39680 66576 39744
rect 66640 39680 66656 39744
rect 66720 39680 66736 39744
rect 66800 39680 66816 39744
rect 66880 39680 66886 39744
rect 66570 39679 66886 39680
rect 5790 39200 6106 39201
rect 5790 39136 5796 39200
rect 5860 39136 5876 39200
rect 5940 39136 5956 39200
rect 6020 39136 6036 39200
rect 6100 39136 6106 39200
rect 5790 39135 6106 39136
rect 36510 39200 36826 39201
rect 36510 39136 36516 39200
rect 36580 39136 36596 39200
rect 36660 39136 36676 39200
rect 36740 39136 36756 39200
rect 36820 39136 36826 39200
rect 36510 39135 36826 39136
rect 67230 39200 67546 39201
rect 67230 39136 67236 39200
rect 67300 39136 67316 39200
rect 67380 39136 67396 39200
rect 67460 39136 67476 39200
rect 67540 39136 67546 39200
rect 67230 39135 67546 39136
rect 77477 38858 77543 38861
rect 79200 38858 80000 38888
rect 77477 38856 80000 38858
rect 77477 38800 77482 38856
rect 77538 38800 80000 38856
rect 77477 38798 80000 38800
rect 77477 38795 77543 38798
rect 79200 38768 80000 38798
rect 5130 38656 5446 38657
rect 5130 38592 5136 38656
rect 5200 38592 5216 38656
rect 5280 38592 5296 38656
rect 5360 38592 5376 38656
rect 5440 38592 5446 38656
rect 5130 38591 5446 38592
rect 35850 38656 36166 38657
rect 35850 38592 35856 38656
rect 35920 38592 35936 38656
rect 36000 38592 36016 38656
rect 36080 38592 36096 38656
rect 36160 38592 36166 38656
rect 35850 38591 36166 38592
rect 66570 38656 66886 38657
rect 66570 38592 66576 38656
rect 66640 38592 66656 38656
rect 66720 38592 66736 38656
rect 66800 38592 66816 38656
rect 66880 38592 66886 38656
rect 66570 38591 66886 38592
rect 77477 38178 77543 38181
rect 79200 38178 80000 38208
rect 77477 38176 80000 38178
rect 77477 38120 77482 38176
rect 77538 38120 80000 38176
rect 77477 38118 80000 38120
rect 77477 38115 77543 38118
rect 5790 38112 6106 38113
rect 5790 38048 5796 38112
rect 5860 38048 5876 38112
rect 5940 38048 5956 38112
rect 6020 38048 6036 38112
rect 6100 38048 6106 38112
rect 5790 38047 6106 38048
rect 36510 38112 36826 38113
rect 36510 38048 36516 38112
rect 36580 38048 36596 38112
rect 36660 38048 36676 38112
rect 36740 38048 36756 38112
rect 36820 38048 36826 38112
rect 36510 38047 36826 38048
rect 67230 38112 67546 38113
rect 67230 38048 67236 38112
rect 67300 38048 67316 38112
rect 67380 38048 67396 38112
rect 67460 38048 67476 38112
rect 67540 38048 67546 38112
rect 79200 38088 80000 38118
rect 67230 38047 67546 38048
rect 5130 37568 5446 37569
rect 5130 37504 5136 37568
rect 5200 37504 5216 37568
rect 5280 37504 5296 37568
rect 5360 37504 5376 37568
rect 5440 37504 5446 37568
rect 5130 37503 5446 37504
rect 35850 37568 36166 37569
rect 35850 37504 35856 37568
rect 35920 37504 35936 37568
rect 36000 37504 36016 37568
rect 36080 37504 36096 37568
rect 36160 37504 36166 37568
rect 35850 37503 36166 37504
rect 66570 37568 66886 37569
rect 66570 37504 66576 37568
rect 66640 37504 66656 37568
rect 66720 37504 66736 37568
rect 66800 37504 66816 37568
rect 66880 37504 66886 37568
rect 66570 37503 66886 37504
rect 77477 37498 77543 37501
rect 79200 37498 80000 37528
rect 77477 37496 80000 37498
rect 77477 37440 77482 37496
rect 77538 37440 80000 37496
rect 77477 37438 80000 37440
rect 77477 37435 77543 37438
rect 79200 37408 80000 37438
rect 5790 37024 6106 37025
rect 5790 36960 5796 37024
rect 5860 36960 5876 37024
rect 5940 36960 5956 37024
rect 6020 36960 6036 37024
rect 6100 36960 6106 37024
rect 5790 36959 6106 36960
rect 36510 37024 36826 37025
rect 36510 36960 36516 37024
rect 36580 36960 36596 37024
rect 36660 36960 36676 37024
rect 36740 36960 36756 37024
rect 36820 36960 36826 37024
rect 36510 36959 36826 36960
rect 67230 37024 67546 37025
rect 67230 36960 67236 37024
rect 67300 36960 67316 37024
rect 67380 36960 67396 37024
rect 67460 36960 67476 37024
rect 67540 36960 67546 37024
rect 67230 36959 67546 36960
rect 77477 36818 77543 36821
rect 79200 36818 80000 36848
rect 77477 36816 80000 36818
rect 77477 36760 77482 36816
rect 77538 36760 80000 36816
rect 77477 36758 80000 36760
rect 77477 36755 77543 36758
rect 79200 36728 80000 36758
rect 5130 36480 5446 36481
rect 5130 36416 5136 36480
rect 5200 36416 5216 36480
rect 5280 36416 5296 36480
rect 5360 36416 5376 36480
rect 5440 36416 5446 36480
rect 5130 36415 5446 36416
rect 35850 36480 36166 36481
rect 35850 36416 35856 36480
rect 35920 36416 35936 36480
rect 36000 36416 36016 36480
rect 36080 36416 36096 36480
rect 36160 36416 36166 36480
rect 35850 36415 36166 36416
rect 66570 36480 66886 36481
rect 66570 36416 66576 36480
rect 66640 36416 66656 36480
rect 66720 36416 66736 36480
rect 66800 36416 66816 36480
rect 66880 36416 66886 36480
rect 66570 36415 66886 36416
rect 5790 35936 6106 35937
rect 5790 35872 5796 35936
rect 5860 35872 5876 35936
rect 5940 35872 5956 35936
rect 6020 35872 6036 35936
rect 6100 35872 6106 35936
rect 5790 35871 6106 35872
rect 36510 35936 36826 35937
rect 36510 35872 36516 35936
rect 36580 35872 36596 35936
rect 36660 35872 36676 35936
rect 36740 35872 36756 35936
rect 36820 35872 36826 35936
rect 36510 35871 36826 35872
rect 67230 35936 67546 35937
rect 67230 35872 67236 35936
rect 67300 35872 67316 35936
rect 67380 35872 67396 35936
rect 67460 35872 67476 35936
rect 67540 35872 67546 35936
rect 67230 35871 67546 35872
rect 0 35458 800 35488
rect 1209 35458 1275 35461
rect 0 35456 1275 35458
rect 0 35400 1214 35456
rect 1270 35400 1275 35456
rect 0 35398 1275 35400
rect 0 35368 800 35398
rect 1209 35395 1275 35398
rect 5130 35392 5446 35393
rect 5130 35328 5136 35392
rect 5200 35328 5216 35392
rect 5280 35328 5296 35392
rect 5360 35328 5376 35392
rect 5440 35328 5446 35392
rect 5130 35327 5446 35328
rect 35850 35392 36166 35393
rect 35850 35328 35856 35392
rect 35920 35328 35936 35392
rect 36000 35328 36016 35392
rect 36080 35328 36096 35392
rect 36160 35328 36166 35392
rect 35850 35327 36166 35328
rect 66570 35392 66886 35393
rect 66570 35328 66576 35392
rect 66640 35328 66656 35392
rect 66720 35328 66736 35392
rect 66800 35328 66816 35392
rect 66880 35328 66886 35392
rect 66570 35327 66886 35328
rect 5790 34848 6106 34849
rect 5790 34784 5796 34848
rect 5860 34784 5876 34848
rect 5940 34784 5956 34848
rect 6020 34784 6036 34848
rect 6100 34784 6106 34848
rect 5790 34783 6106 34784
rect 36510 34848 36826 34849
rect 36510 34784 36516 34848
rect 36580 34784 36596 34848
rect 36660 34784 36676 34848
rect 36740 34784 36756 34848
rect 36820 34784 36826 34848
rect 36510 34783 36826 34784
rect 67230 34848 67546 34849
rect 67230 34784 67236 34848
rect 67300 34784 67316 34848
rect 67380 34784 67396 34848
rect 67460 34784 67476 34848
rect 67540 34784 67546 34848
rect 67230 34783 67546 34784
rect 5130 34304 5446 34305
rect 5130 34240 5136 34304
rect 5200 34240 5216 34304
rect 5280 34240 5296 34304
rect 5360 34240 5376 34304
rect 5440 34240 5446 34304
rect 5130 34239 5446 34240
rect 35850 34304 36166 34305
rect 35850 34240 35856 34304
rect 35920 34240 35936 34304
rect 36000 34240 36016 34304
rect 36080 34240 36096 34304
rect 36160 34240 36166 34304
rect 35850 34239 36166 34240
rect 66570 34304 66886 34305
rect 66570 34240 66576 34304
rect 66640 34240 66656 34304
rect 66720 34240 66736 34304
rect 66800 34240 66816 34304
rect 66880 34240 66886 34304
rect 66570 34239 66886 34240
rect 77477 34098 77543 34101
rect 79200 34098 80000 34128
rect 77477 34096 80000 34098
rect 77477 34040 77482 34096
rect 77538 34040 80000 34096
rect 77477 34038 80000 34040
rect 77477 34035 77543 34038
rect 79200 34008 80000 34038
rect 5790 33760 6106 33761
rect 5790 33696 5796 33760
rect 5860 33696 5876 33760
rect 5940 33696 5956 33760
rect 6020 33696 6036 33760
rect 6100 33696 6106 33760
rect 5790 33695 6106 33696
rect 36510 33760 36826 33761
rect 36510 33696 36516 33760
rect 36580 33696 36596 33760
rect 36660 33696 36676 33760
rect 36740 33696 36756 33760
rect 36820 33696 36826 33760
rect 36510 33695 36826 33696
rect 67230 33760 67546 33761
rect 67230 33696 67236 33760
rect 67300 33696 67316 33760
rect 67380 33696 67396 33760
rect 67460 33696 67476 33760
rect 67540 33696 67546 33760
rect 67230 33695 67546 33696
rect 5130 33216 5446 33217
rect 5130 33152 5136 33216
rect 5200 33152 5216 33216
rect 5280 33152 5296 33216
rect 5360 33152 5376 33216
rect 5440 33152 5446 33216
rect 5130 33151 5446 33152
rect 35850 33216 36166 33217
rect 35850 33152 35856 33216
rect 35920 33152 35936 33216
rect 36000 33152 36016 33216
rect 36080 33152 36096 33216
rect 36160 33152 36166 33216
rect 35850 33151 36166 33152
rect 66570 33216 66886 33217
rect 66570 33152 66576 33216
rect 66640 33152 66656 33216
rect 66720 33152 66736 33216
rect 66800 33152 66816 33216
rect 66880 33152 66886 33216
rect 66570 33151 66886 33152
rect 5790 32672 6106 32673
rect 5790 32608 5796 32672
rect 5860 32608 5876 32672
rect 5940 32608 5956 32672
rect 6020 32608 6036 32672
rect 6100 32608 6106 32672
rect 5790 32607 6106 32608
rect 36510 32672 36826 32673
rect 36510 32608 36516 32672
rect 36580 32608 36596 32672
rect 36660 32608 36676 32672
rect 36740 32608 36756 32672
rect 36820 32608 36826 32672
rect 36510 32607 36826 32608
rect 67230 32672 67546 32673
rect 67230 32608 67236 32672
rect 67300 32608 67316 32672
rect 67380 32608 67396 32672
rect 67460 32608 67476 32672
rect 67540 32608 67546 32672
rect 67230 32607 67546 32608
rect 5130 32128 5446 32129
rect 0 32058 800 32088
rect 5130 32064 5136 32128
rect 5200 32064 5216 32128
rect 5280 32064 5296 32128
rect 5360 32064 5376 32128
rect 5440 32064 5446 32128
rect 5130 32063 5446 32064
rect 35850 32128 36166 32129
rect 35850 32064 35856 32128
rect 35920 32064 35936 32128
rect 36000 32064 36016 32128
rect 36080 32064 36096 32128
rect 36160 32064 36166 32128
rect 35850 32063 36166 32064
rect 66570 32128 66886 32129
rect 66570 32064 66576 32128
rect 66640 32064 66656 32128
rect 66720 32064 66736 32128
rect 66800 32064 66816 32128
rect 66880 32064 66886 32128
rect 66570 32063 66886 32064
rect 1209 32058 1275 32061
rect 0 32056 1275 32058
rect 0 32000 1214 32056
rect 1270 32000 1275 32056
rect 0 31998 1275 32000
rect 0 31968 800 31998
rect 1209 31995 1275 31998
rect 5790 31584 6106 31585
rect 5790 31520 5796 31584
rect 5860 31520 5876 31584
rect 5940 31520 5956 31584
rect 6020 31520 6036 31584
rect 6100 31520 6106 31584
rect 5790 31519 6106 31520
rect 36510 31584 36826 31585
rect 36510 31520 36516 31584
rect 36580 31520 36596 31584
rect 36660 31520 36676 31584
rect 36740 31520 36756 31584
rect 36820 31520 36826 31584
rect 36510 31519 36826 31520
rect 67230 31584 67546 31585
rect 67230 31520 67236 31584
rect 67300 31520 67316 31584
rect 67380 31520 67396 31584
rect 67460 31520 67476 31584
rect 67540 31520 67546 31584
rect 67230 31519 67546 31520
rect 5130 31040 5446 31041
rect 5130 30976 5136 31040
rect 5200 30976 5216 31040
rect 5280 30976 5296 31040
rect 5360 30976 5376 31040
rect 5440 30976 5446 31040
rect 5130 30975 5446 30976
rect 35850 31040 36166 31041
rect 35850 30976 35856 31040
rect 35920 30976 35936 31040
rect 36000 30976 36016 31040
rect 36080 30976 36096 31040
rect 36160 30976 36166 31040
rect 35850 30975 36166 30976
rect 66570 31040 66886 31041
rect 66570 30976 66576 31040
rect 66640 30976 66656 31040
rect 66720 30976 66736 31040
rect 66800 30976 66816 31040
rect 66880 30976 66886 31040
rect 66570 30975 66886 30976
rect 5790 30496 6106 30497
rect 5790 30432 5796 30496
rect 5860 30432 5876 30496
rect 5940 30432 5956 30496
rect 6020 30432 6036 30496
rect 6100 30432 6106 30496
rect 5790 30431 6106 30432
rect 36510 30496 36826 30497
rect 36510 30432 36516 30496
rect 36580 30432 36596 30496
rect 36660 30432 36676 30496
rect 36740 30432 36756 30496
rect 36820 30432 36826 30496
rect 36510 30431 36826 30432
rect 67230 30496 67546 30497
rect 67230 30432 67236 30496
rect 67300 30432 67316 30496
rect 67380 30432 67396 30496
rect 67460 30432 67476 30496
rect 67540 30432 67546 30496
rect 67230 30431 67546 30432
rect 5130 29952 5446 29953
rect 5130 29888 5136 29952
rect 5200 29888 5216 29952
rect 5280 29888 5296 29952
rect 5360 29888 5376 29952
rect 5440 29888 5446 29952
rect 5130 29887 5446 29888
rect 35850 29952 36166 29953
rect 35850 29888 35856 29952
rect 35920 29888 35936 29952
rect 36000 29888 36016 29952
rect 36080 29888 36096 29952
rect 36160 29888 36166 29952
rect 35850 29887 36166 29888
rect 66570 29952 66886 29953
rect 66570 29888 66576 29952
rect 66640 29888 66656 29952
rect 66720 29888 66736 29952
rect 66800 29888 66816 29952
rect 66880 29888 66886 29952
rect 66570 29887 66886 29888
rect 5790 29408 6106 29409
rect 5790 29344 5796 29408
rect 5860 29344 5876 29408
rect 5940 29344 5956 29408
rect 6020 29344 6036 29408
rect 6100 29344 6106 29408
rect 5790 29343 6106 29344
rect 36510 29408 36826 29409
rect 36510 29344 36516 29408
rect 36580 29344 36596 29408
rect 36660 29344 36676 29408
rect 36740 29344 36756 29408
rect 36820 29344 36826 29408
rect 36510 29343 36826 29344
rect 67230 29408 67546 29409
rect 67230 29344 67236 29408
rect 67300 29344 67316 29408
rect 67380 29344 67396 29408
rect 67460 29344 67476 29408
rect 67540 29344 67546 29408
rect 67230 29343 67546 29344
rect 5130 28864 5446 28865
rect 5130 28800 5136 28864
rect 5200 28800 5216 28864
rect 5280 28800 5296 28864
rect 5360 28800 5376 28864
rect 5440 28800 5446 28864
rect 5130 28799 5446 28800
rect 35850 28864 36166 28865
rect 35850 28800 35856 28864
rect 35920 28800 35936 28864
rect 36000 28800 36016 28864
rect 36080 28800 36096 28864
rect 36160 28800 36166 28864
rect 35850 28799 36166 28800
rect 66570 28864 66886 28865
rect 66570 28800 66576 28864
rect 66640 28800 66656 28864
rect 66720 28800 66736 28864
rect 66800 28800 66816 28864
rect 66880 28800 66886 28864
rect 66570 28799 66886 28800
rect 0 28658 800 28688
rect 2313 28658 2379 28661
rect 0 28656 2379 28658
rect 0 28600 2318 28656
rect 2374 28600 2379 28656
rect 0 28598 2379 28600
rect 0 28568 800 28598
rect 2313 28595 2379 28598
rect 5790 28320 6106 28321
rect 5790 28256 5796 28320
rect 5860 28256 5876 28320
rect 5940 28256 5956 28320
rect 6020 28256 6036 28320
rect 6100 28256 6106 28320
rect 5790 28255 6106 28256
rect 36510 28320 36826 28321
rect 36510 28256 36516 28320
rect 36580 28256 36596 28320
rect 36660 28256 36676 28320
rect 36740 28256 36756 28320
rect 36820 28256 36826 28320
rect 36510 28255 36826 28256
rect 67230 28320 67546 28321
rect 67230 28256 67236 28320
rect 67300 28256 67316 28320
rect 67380 28256 67396 28320
rect 67460 28256 67476 28320
rect 67540 28256 67546 28320
rect 67230 28255 67546 28256
rect 0 27978 800 28008
rect 1209 27978 1275 27981
rect 0 27976 1275 27978
rect 0 27920 1214 27976
rect 1270 27920 1275 27976
rect 0 27918 1275 27920
rect 0 27888 800 27918
rect 1209 27915 1275 27918
rect 5130 27776 5446 27777
rect 5130 27712 5136 27776
rect 5200 27712 5216 27776
rect 5280 27712 5296 27776
rect 5360 27712 5376 27776
rect 5440 27712 5446 27776
rect 5130 27711 5446 27712
rect 35850 27776 36166 27777
rect 35850 27712 35856 27776
rect 35920 27712 35936 27776
rect 36000 27712 36016 27776
rect 36080 27712 36096 27776
rect 36160 27712 36166 27776
rect 35850 27711 36166 27712
rect 66570 27776 66886 27777
rect 66570 27712 66576 27776
rect 66640 27712 66656 27776
rect 66720 27712 66736 27776
rect 66800 27712 66816 27776
rect 66880 27712 66886 27776
rect 66570 27711 66886 27712
rect 5790 27232 6106 27233
rect 5790 27168 5796 27232
rect 5860 27168 5876 27232
rect 5940 27168 5956 27232
rect 6020 27168 6036 27232
rect 6100 27168 6106 27232
rect 5790 27167 6106 27168
rect 36510 27232 36826 27233
rect 36510 27168 36516 27232
rect 36580 27168 36596 27232
rect 36660 27168 36676 27232
rect 36740 27168 36756 27232
rect 36820 27168 36826 27232
rect 36510 27167 36826 27168
rect 67230 27232 67546 27233
rect 67230 27168 67236 27232
rect 67300 27168 67316 27232
rect 67380 27168 67396 27232
rect 67460 27168 67476 27232
rect 67540 27168 67546 27232
rect 67230 27167 67546 27168
rect 5130 26688 5446 26689
rect 0 26618 800 26648
rect 5130 26624 5136 26688
rect 5200 26624 5216 26688
rect 5280 26624 5296 26688
rect 5360 26624 5376 26688
rect 5440 26624 5446 26688
rect 5130 26623 5446 26624
rect 35850 26688 36166 26689
rect 35850 26624 35856 26688
rect 35920 26624 35936 26688
rect 36000 26624 36016 26688
rect 36080 26624 36096 26688
rect 36160 26624 36166 26688
rect 35850 26623 36166 26624
rect 66570 26688 66886 26689
rect 66570 26624 66576 26688
rect 66640 26624 66656 26688
rect 66720 26624 66736 26688
rect 66800 26624 66816 26688
rect 66880 26624 66886 26688
rect 66570 26623 66886 26624
rect 1209 26618 1275 26621
rect 0 26616 1275 26618
rect 0 26560 1214 26616
rect 1270 26560 1275 26616
rect 0 26558 1275 26560
rect 0 26528 800 26558
rect 1209 26555 1275 26558
rect 5790 26144 6106 26145
rect 5790 26080 5796 26144
rect 5860 26080 5876 26144
rect 5940 26080 5956 26144
rect 6020 26080 6036 26144
rect 6100 26080 6106 26144
rect 5790 26079 6106 26080
rect 36510 26144 36826 26145
rect 36510 26080 36516 26144
rect 36580 26080 36596 26144
rect 36660 26080 36676 26144
rect 36740 26080 36756 26144
rect 36820 26080 36826 26144
rect 36510 26079 36826 26080
rect 67230 26144 67546 26145
rect 67230 26080 67236 26144
rect 67300 26080 67316 26144
rect 67380 26080 67396 26144
rect 67460 26080 67476 26144
rect 67540 26080 67546 26144
rect 67230 26079 67546 26080
rect 0 25938 800 25968
rect 2313 25938 2379 25941
rect 0 25936 2379 25938
rect 0 25880 2318 25936
rect 2374 25880 2379 25936
rect 0 25878 2379 25880
rect 0 25848 800 25878
rect 2313 25875 2379 25878
rect 5130 25600 5446 25601
rect 5130 25536 5136 25600
rect 5200 25536 5216 25600
rect 5280 25536 5296 25600
rect 5360 25536 5376 25600
rect 5440 25536 5446 25600
rect 5130 25535 5446 25536
rect 35850 25600 36166 25601
rect 35850 25536 35856 25600
rect 35920 25536 35936 25600
rect 36000 25536 36016 25600
rect 36080 25536 36096 25600
rect 36160 25536 36166 25600
rect 35850 25535 36166 25536
rect 66570 25600 66886 25601
rect 66570 25536 66576 25600
rect 66640 25536 66656 25600
rect 66720 25536 66736 25600
rect 66800 25536 66816 25600
rect 66880 25536 66886 25600
rect 66570 25535 66886 25536
rect 5790 25056 6106 25057
rect 5790 24992 5796 25056
rect 5860 24992 5876 25056
rect 5940 24992 5956 25056
rect 6020 24992 6036 25056
rect 6100 24992 6106 25056
rect 5790 24991 6106 24992
rect 36510 25056 36826 25057
rect 36510 24992 36516 25056
rect 36580 24992 36596 25056
rect 36660 24992 36676 25056
rect 36740 24992 36756 25056
rect 36820 24992 36826 25056
rect 36510 24991 36826 24992
rect 67230 25056 67546 25057
rect 67230 24992 67236 25056
rect 67300 24992 67316 25056
rect 67380 24992 67396 25056
rect 67460 24992 67476 25056
rect 67540 24992 67546 25056
rect 67230 24991 67546 24992
rect 5130 24512 5446 24513
rect 5130 24448 5136 24512
rect 5200 24448 5216 24512
rect 5280 24448 5296 24512
rect 5360 24448 5376 24512
rect 5440 24448 5446 24512
rect 5130 24447 5446 24448
rect 35850 24512 36166 24513
rect 35850 24448 35856 24512
rect 35920 24448 35936 24512
rect 36000 24448 36016 24512
rect 36080 24448 36096 24512
rect 36160 24448 36166 24512
rect 35850 24447 36166 24448
rect 66570 24512 66886 24513
rect 66570 24448 66576 24512
rect 66640 24448 66656 24512
rect 66720 24448 66736 24512
rect 66800 24448 66816 24512
rect 66880 24448 66886 24512
rect 66570 24447 66886 24448
rect 5790 23968 6106 23969
rect 5790 23904 5796 23968
rect 5860 23904 5876 23968
rect 5940 23904 5956 23968
rect 6020 23904 6036 23968
rect 6100 23904 6106 23968
rect 5790 23903 6106 23904
rect 36510 23968 36826 23969
rect 36510 23904 36516 23968
rect 36580 23904 36596 23968
rect 36660 23904 36676 23968
rect 36740 23904 36756 23968
rect 36820 23904 36826 23968
rect 36510 23903 36826 23904
rect 67230 23968 67546 23969
rect 67230 23904 67236 23968
rect 67300 23904 67316 23968
rect 67380 23904 67396 23968
rect 67460 23904 67476 23968
rect 67540 23904 67546 23968
rect 67230 23903 67546 23904
rect 5130 23424 5446 23425
rect 5130 23360 5136 23424
rect 5200 23360 5216 23424
rect 5280 23360 5296 23424
rect 5360 23360 5376 23424
rect 5440 23360 5446 23424
rect 5130 23359 5446 23360
rect 35850 23424 36166 23425
rect 35850 23360 35856 23424
rect 35920 23360 35936 23424
rect 36000 23360 36016 23424
rect 36080 23360 36096 23424
rect 36160 23360 36166 23424
rect 35850 23359 36166 23360
rect 66570 23424 66886 23425
rect 66570 23360 66576 23424
rect 66640 23360 66656 23424
rect 66720 23360 66736 23424
rect 66800 23360 66816 23424
rect 66880 23360 66886 23424
rect 66570 23359 66886 23360
rect 0 23218 800 23248
rect 2313 23218 2379 23221
rect 0 23216 2379 23218
rect 0 23160 2318 23216
rect 2374 23160 2379 23216
rect 0 23158 2379 23160
rect 0 23128 800 23158
rect 2313 23155 2379 23158
rect 5790 22880 6106 22881
rect 5790 22816 5796 22880
rect 5860 22816 5876 22880
rect 5940 22816 5956 22880
rect 6020 22816 6036 22880
rect 6100 22816 6106 22880
rect 5790 22815 6106 22816
rect 36510 22880 36826 22881
rect 36510 22816 36516 22880
rect 36580 22816 36596 22880
rect 36660 22816 36676 22880
rect 36740 22816 36756 22880
rect 36820 22816 36826 22880
rect 36510 22815 36826 22816
rect 67230 22880 67546 22881
rect 67230 22816 67236 22880
rect 67300 22816 67316 22880
rect 67380 22816 67396 22880
rect 67460 22816 67476 22880
rect 67540 22816 67546 22880
rect 67230 22815 67546 22816
rect 5130 22336 5446 22337
rect 5130 22272 5136 22336
rect 5200 22272 5216 22336
rect 5280 22272 5296 22336
rect 5360 22272 5376 22336
rect 5440 22272 5446 22336
rect 5130 22271 5446 22272
rect 35850 22336 36166 22337
rect 35850 22272 35856 22336
rect 35920 22272 35936 22336
rect 36000 22272 36016 22336
rect 36080 22272 36096 22336
rect 36160 22272 36166 22336
rect 35850 22271 36166 22272
rect 66570 22336 66886 22337
rect 66570 22272 66576 22336
rect 66640 22272 66656 22336
rect 66720 22272 66736 22336
rect 66800 22272 66816 22336
rect 66880 22272 66886 22336
rect 66570 22271 66886 22272
rect 5790 21792 6106 21793
rect 5790 21728 5796 21792
rect 5860 21728 5876 21792
rect 5940 21728 5956 21792
rect 6020 21728 6036 21792
rect 6100 21728 6106 21792
rect 5790 21727 6106 21728
rect 36510 21792 36826 21793
rect 36510 21728 36516 21792
rect 36580 21728 36596 21792
rect 36660 21728 36676 21792
rect 36740 21728 36756 21792
rect 36820 21728 36826 21792
rect 36510 21727 36826 21728
rect 67230 21792 67546 21793
rect 67230 21728 67236 21792
rect 67300 21728 67316 21792
rect 67380 21728 67396 21792
rect 67460 21728 67476 21792
rect 67540 21728 67546 21792
rect 67230 21727 67546 21728
rect 5130 21248 5446 21249
rect 5130 21184 5136 21248
rect 5200 21184 5216 21248
rect 5280 21184 5296 21248
rect 5360 21184 5376 21248
rect 5440 21184 5446 21248
rect 5130 21183 5446 21184
rect 35850 21248 36166 21249
rect 35850 21184 35856 21248
rect 35920 21184 35936 21248
rect 36000 21184 36016 21248
rect 36080 21184 36096 21248
rect 36160 21184 36166 21248
rect 35850 21183 36166 21184
rect 66570 21248 66886 21249
rect 66570 21184 66576 21248
rect 66640 21184 66656 21248
rect 66720 21184 66736 21248
rect 66800 21184 66816 21248
rect 66880 21184 66886 21248
rect 66570 21183 66886 21184
rect 77569 21178 77635 21181
rect 79200 21178 80000 21208
rect 77569 21176 80000 21178
rect 77569 21120 77574 21176
rect 77630 21120 80000 21176
rect 77569 21118 80000 21120
rect 77569 21115 77635 21118
rect 79200 21088 80000 21118
rect 5790 20704 6106 20705
rect 5790 20640 5796 20704
rect 5860 20640 5876 20704
rect 5940 20640 5956 20704
rect 6020 20640 6036 20704
rect 6100 20640 6106 20704
rect 5790 20639 6106 20640
rect 36510 20704 36826 20705
rect 36510 20640 36516 20704
rect 36580 20640 36596 20704
rect 36660 20640 36676 20704
rect 36740 20640 36756 20704
rect 36820 20640 36826 20704
rect 36510 20639 36826 20640
rect 67230 20704 67546 20705
rect 67230 20640 67236 20704
rect 67300 20640 67316 20704
rect 67380 20640 67396 20704
rect 67460 20640 67476 20704
rect 67540 20640 67546 20704
rect 67230 20639 67546 20640
rect 5130 20160 5446 20161
rect 5130 20096 5136 20160
rect 5200 20096 5216 20160
rect 5280 20096 5296 20160
rect 5360 20096 5376 20160
rect 5440 20096 5446 20160
rect 5130 20095 5446 20096
rect 35850 20160 36166 20161
rect 35850 20096 35856 20160
rect 35920 20096 35936 20160
rect 36000 20096 36016 20160
rect 36080 20096 36096 20160
rect 36160 20096 36166 20160
rect 35850 20095 36166 20096
rect 66570 20160 66886 20161
rect 66570 20096 66576 20160
rect 66640 20096 66656 20160
rect 66720 20096 66736 20160
rect 66800 20096 66816 20160
rect 66880 20096 66886 20160
rect 66570 20095 66886 20096
rect 5790 19616 6106 19617
rect 5790 19552 5796 19616
rect 5860 19552 5876 19616
rect 5940 19552 5956 19616
rect 6020 19552 6036 19616
rect 6100 19552 6106 19616
rect 5790 19551 6106 19552
rect 36510 19616 36826 19617
rect 36510 19552 36516 19616
rect 36580 19552 36596 19616
rect 36660 19552 36676 19616
rect 36740 19552 36756 19616
rect 36820 19552 36826 19616
rect 36510 19551 36826 19552
rect 67230 19616 67546 19617
rect 67230 19552 67236 19616
rect 67300 19552 67316 19616
rect 67380 19552 67396 19616
rect 67460 19552 67476 19616
rect 67540 19552 67546 19616
rect 67230 19551 67546 19552
rect 5130 19072 5446 19073
rect 5130 19008 5136 19072
rect 5200 19008 5216 19072
rect 5280 19008 5296 19072
rect 5360 19008 5376 19072
rect 5440 19008 5446 19072
rect 5130 19007 5446 19008
rect 35850 19072 36166 19073
rect 35850 19008 35856 19072
rect 35920 19008 35936 19072
rect 36000 19008 36016 19072
rect 36080 19008 36096 19072
rect 36160 19008 36166 19072
rect 35850 19007 36166 19008
rect 66570 19072 66886 19073
rect 66570 19008 66576 19072
rect 66640 19008 66656 19072
rect 66720 19008 66736 19072
rect 66800 19008 66816 19072
rect 66880 19008 66886 19072
rect 66570 19007 66886 19008
rect 5790 18528 6106 18529
rect 5790 18464 5796 18528
rect 5860 18464 5876 18528
rect 5940 18464 5956 18528
rect 6020 18464 6036 18528
rect 6100 18464 6106 18528
rect 5790 18463 6106 18464
rect 36510 18528 36826 18529
rect 36510 18464 36516 18528
rect 36580 18464 36596 18528
rect 36660 18464 36676 18528
rect 36740 18464 36756 18528
rect 36820 18464 36826 18528
rect 36510 18463 36826 18464
rect 67230 18528 67546 18529
rect 67230 18464 67236 18528
rect 67300 18464 67316 18528
rect 67380 18464 67396 18528
rect 67460 18464 67476 18528
rect 67540 18464 67546 18528
rect 67230 18463 67546 18464
rect 5130 17984 5446 17985
rect 5130 17920 5136 17984
rect 5200 17920 5216 17984
rect 5280 17920 5296 17984
rect 5360 17920 5376 17984
rect 5440 17920 5446 17984
rect 5130 17919 5446 17920
rect 35850 17984 36166 17985
rect 35850 17920 35856 17984
rect 35920 17920 35936 17984
rect 36000 17920 36016 17984
rect 36080 17920 36096 17984
rect 36160 17920 36166 17984
rect 35850 17919 36166 17920
rect 66570 17984 66886 17985
rect 66570 17920 66576 17984
rect 66640 17920 66656 17984
rect 66720 17920 66736 17984
rect 66800 17920 66816 17984
rect 66880 17920 66886 17984
rect 66570 17919 66886 17920
rect 5790 17440 6106 17441
rect 5790 17376 5796 17440
rect 5860 17376 5876 17440
rect 5940 17376 5956 17440
rect 6020 17376 6036 17440
rect 6100 17376 6106 17440
rect 5790 17375 6106 17376
rect 36510 17440 36826 17441
rect 36510 17376 36516 17440
rect 36580 17376 36596 17440
rect 36660 17376 36676 17440
rect 36740 17376 36756 17440
rect 36820 17376 36826 17440
rect 36510 17375 36826 17376
rect 67230 17440 67546 17441
rect 67230 17376 67236 17440
rect 67300 17376 67316 17440
rect 67380 17376 67396 17440
rect 67460 17376 67476 17440
rect 67540 17376 67546 17440
rect 67230 17375 67546 17376
rect 5130 16896 5446 16897
rect 5130 16832 5136 16896
rect 5200 16832 5216 16896
rect 5280 16832 5296 16896
rect 5360 16832 5376 16896
rect 5440 16832 5446 16896
rect 5130 16831 5446 16832
rect 35850 16896 36166 16897
rect 35850 16832 35856 16896
rect 35920 16832 35936 16896
rect 36000 16832 36016 16896
rect 36080 16832 36096 16896
rect 36160 16832 36166 16896
rect 35850 16831 36166 16832
rect 66570 16896 66886 16897
rect 66570 16832 66576 16896
rect 66640 16832 66656 16896
rect 66720 16832 66736 16896
rect 66800 16832 66816 16896
rect 66880 16832 66886 16896
rect 66570 16831 66886 16832
rect 77569 16418 77635 16421
rect 79200 16418 80000 16448
rect 77569 16416 80000 16418
rect 77569 16360 77574 16416
rect 77630 16360 80000 16416
rect 77569 16358 80000 16360
rect 77569 16355 77635 16358
rect 5790 16352 6106 16353
rect 5790 16288 5796 16352
rect 5860 16288 5876 16352
rect 5940 16288 5956 16352
rect 6020 16288 6036 16352
rect 6100 16288 6106 16352
rect 5790 16287 6106 16288
rect 36510 16352 36826 16353
rect 36510 16288 36516 16352
rect 36580 16288 36596 16352
rect 36660 16288 36676 16352
rect 36740 16288 36756 16352
rect 36820 16288 36826 16352
rect 36510 16287 36826 16288
rect 67230 16352 67546 16353
rect 67230 16288 67236 16352
rect 67300 16288 67316 16352
rect 67380 16288 67396 16352
rect 67460 16288 67476 16352
rect 67540 16288 67546 16352
rect 79200 16328 80000 16358
rect 67230 16287 67546 16288
rect 5130 15808 5446 15809
rect 5130 15744 5136 15808
rect 5200 15744 5216 15808
rect 5280 15744 5296 15808
rect 5360 15744 5376 15808
rect 5440 15744 5446 15808
rect 5130 15743 5446 15744
rect 35850 15808 36166 15809
rect 35850 15744 35856 15808
rect 35920 15744 35936 15808
rect 36000 15744 36016 15808
rect 36080 15744 36096 15808
rect 36160 15744 36166 15808
rect 35850 15743 36166 15744
rect 66570 15808 66886 15809
rect 66570 15744 66576 15808
rect 66640 15744 66656 15808
rect 66720 15744 66736 15808
rect 66800 15744 66816 15808
rect 66880 15744 66886 15808
rect 66570 15743 66886 15744
rect 5790 15264 6106 15265
rect 5790 15200 5796 15264
rect 5860 15200 5876 15264
rect 5940 15200 5956 15264
rect 6020 15200 6036 15264
rect 6100 15200 6106 15264
rect 5790 15199 6106 15200
rect 36510 15264 36826 15265
rect 36510 15200 36516 15264
rect 36580 15200 36596 15264
rect 36660 15200 36676 15264
rect 36740 15200 36756 15264
rect 36820 15200 36826 15264
rect 36510 15199 36826 15200
rect 67230 15264 67546 15265
rect 67230 15200 67236 15264
rect 67300 15200 67316 15264
rect 67380 15200 67396 15264
rect 67460 15200 67476 15264
rect 67540 15200 67546 15264
rect 67230 15199 67546 15200
rect 5130 14720 5446 14721
rect 5130 14656 5136 14720
rect 5200 14656 5216 14720
rect 5280 14656 5296 14720
rect 5360 14656 5376 14720
rect 5440 14656 5446 14720
rect 5130 14655 5446 14656
rect 35850 14720 36166 14721
rect 35850 14656 35856 14720
rect 35920 14656 35936 14720
rect 36000 14656 36016 14720
rect 36080 14656 36096 14720
rect 36160 14656 36166 14720
rect 35850 14655 36166 14656
rect 66570 14720 66886 14721
rect 66570 14656 66576 14720
rect 66640 14656 66656 14720
rect 66720 14656 66736 14720
rect 66800 14656 66816 14720
rect 66880 14656 66886 14720
rect 66570 14655 66886 14656
rect 5790 14176 6106 14177
rect 5790 14112 5796 14176
rect 5860 14112 5876 14176
rect 5940 14112 5956 14176
rect 6020 14112 6036 14176
rect 6100 14112 6106 14176
rect 5790 14111 6106 14112
rect 36510 14176 36826 14177
rect 36510 14112 36516 14176
rect 36580 14112 36596 14176
rect 36660 14112 36676 14176
rect 36740 14112 36756 14176
rect 36820 14112 36826 14176
rect 36510 14111 36826 14112
rect 67230 14176 67546 14177
rect 67230 14112 67236 14176
rect 67300 14112 67316 14176
rect 67380 14112 67396 14176
rect 67460 14112 67476 14176
rect 67540 14112 67546 14176
rect 67230 14111 67546 14112
rect 5130 13632 5446 13633
rect 5130 13568 5136 13632
rect 5200 13568 5216 13632
rect 5280 13568 5296 13632
rect 5360 13568 5376 13632
rect 5440 13568 5446 13632
rect 5130 13567 5446 13568
rect 35850 13632 36166 13633
rect 35850 13568 35856 13632
rect 35920 13568 35936 13632
rect 36000 13568 36016 13632
rect 36080 13568 36096 13632
rect 36160 13568 36166 13632
rect 35850 13567 36166 13568
rect 66570 13632 66886 13633
rect 66570 13568 66576 13632
rect 66640 13568 66656 13632
rect 66720 13568 66736 13632
rect 66800 13568 66816 13632
rect 66880 13568 66886 13632
rect 66570 13567 66886 13568
rect 5790 13088 6106 13089
rect 5790 13024 5796 13088
rect 5860 13024 5876 13088
rect 5940 13024 5956 13088
rect 6020 13024 6036 13088
rect 6100 13024 6106 13088
rect 5790 13023 6106 13024
rect 36510 13088 36826 13089
rect 36510 13024 36516 13088
rect 36580 13024 36596 13088
rect 36660 13024 36676 13088
rect 36740 13024 36756 13088
rect 36820 13024 36826 13088
rect 36510 13023 36826 13024
rect 67230 13088 67546 13089
rect 67230 13024 67236 13088
rect 67300 13024 67316 13088
rect 67380 13024 67396 13088
rect 67460 13024 67476 13088
rect 67540 13024 67546 13088
rect 67230 13023 67546 13024
rect 5130 12544 5446 12545
rect 5130 12480 5136 12544
rect 5200 12480 5216 12544
rect 5280 12480 5296 12544
rect 5360 12480 5376 12544
rect 5440 12480 5446 12544
rect 5130 12479 5446 12480
rect 35850 12544 36166 12545
rect 35850 12480 35856 12544
rect 35920 12480 35936 12544
rect 36000 12480 36016 12544
rect 36080 12480 36096 12544
rect 36160 12480 36166 12544
rect 35850 12479 36166 12480
rect 66570 12544 66886 12545
rect 66570 12480 66576 12544
rect 66640 12480 66656 12544
rect 66720 12480 66736 12544
rect 66800 12480 66816 12544
rect 66880 12480 66886 12544
rect 66570 12479 66886 12480
rect 5790 12000 6106 12001
rect 5790 11936 5796 12000
rect 5860 11936 5876 12000
rect 5940 11936 5956 12000
rect 6020 11936 6036 12000
rect 6100 11936 6106 12000
rect 5790 11935 6106 11936
rect 36510 12000 36826 12001
rect 36510 11936 36516 12000
rect 36580 11936 36596 12000
rect 36660 11936 36676 12000
rect 36740 11936 36756 12000
rect 36820 11936 36826 12000
rect 36510 11935 36826 11936
rect 67230 12000 67546 12001
rect 67230 11936 67236 12000
rect 67300 11936 67316 12000
rect 67380 11936 67396 12000
rect 67460 11936 67476 12000
rect 67540 11936 67546 12000
rect 67230 11935 67546 11936
rect 5130 11456 5446 11457
rect 5130 11392 5136 11456
rect 5200 11392 5216 11456
rect 5280 11392 5296 11456
rect 5360 11392 5376 11456
rect 5440 11392 5446 11456
rect 5130 11391 5446 11392
rect 35850 11456 36166 11457
rect 35850 11392 35856 11456
rect 35920 11392 35936 11456
rect 36000 11392 36016 11456
rect 36080 11392 36096 11456
rect 36160 11392 36166 11456
rect 35850 11391 36166 11392
rect 66570 11456 66886 11457
rect 66570 11392 66576 11456
rect 66640 11392 66656 11456
rect 66720 11392 66736 11456
rect 66800 11392 66816 11456
rect 66880 11392 66886 11456
rect 66570 11391 66886 11392
rect 5790 10912 6106 10913
rect 5790 10848 5796 10912
rect 5860 10848 5876 10912
rect 5940 10848 5956 10912
rect 6020 10848 6036 10912
rect 6100 10848 6106 10912
rect 5790 10847 6106 10848
rect 36510 10912 36826 10913
rect 36510 10848 36516 10912
rect 36580 10848 36596 10912
rect 36660 10848 36676 10912
rect 36740 10848 36756 10912
rect 36820 10848 36826 10912
rect 36510 10847 36826 10848
rect 67230 10912 67546 10913
rect 67230 10848 67236 10912
rect 67300 10848 67316 10912
rect 67380 10848 67396 10912
rect 67460 10848 67476 10912
rect 67540 10848 67546 10912
rect 67230 10847 67546 10848
rect 5130 10368 5446 10369
rect 5130 10304 5136 10368
rect 5200 10304 5216 10368
rect 5280 10304 5296 10368
rect 5360 10304 5376 10368
rect 5440 10304 5446 10368
rect 5130 10303 5446 10304
rect 35850 10368 36166 10369
rect 35850 10304 35856 10368
rect 35920 10304 35936 10368
rect 36000 10304 36016 10368
rect 36080 10304 36096 10368
rect 36160 10304 36166 10368
rect 35850 10303 36166 10304
rect 66570 10368 66886 10369
rect 66570 10304 66576 10368
rect 66640 10304 66656 10368
rect 66720 10304 66736 10368
rect 66800 10304 66816 10368
rect 66880 10304 66886 10368
rect 66570 10303 66886 10304
rect 5790 9824 6106 9825
rect 5790 9760 5796 9824
rect 5860 9760 5876 9824
rect 5940 9760 5956 9824
rect 6020 9760 6036 9824
rect 6100 9760 6106 9824
rect 5790 9759 6106 9760
rect 36510 9824 36826 9825
rect 36510 9760 36516 9824
rect 36580 9760 36596 9824
rect 36660 9760 36676 9824
rect 36740 9760 36756 9824
rect 36820 9760 36826 9824
rect 36510 9759 36826 9760
rect 67230 9824 67546 9825
rect 67230 9760 67236 9824
rect 67300 9760 67316 9824
rect 67380 9760 67396 9824
rect 67460 9760 67476 9824
rect 67540 9760 67546 9824
rect 67230 9759 67546 9760
rect 5130 9280 5446 9281
rect 5130 9216 5136 9280
rect 5200 9216 5216 9280
rect 5280 9216 5296 9280
rect 5360 9216 5376 9280
rect 5440 9216 5446 9280
rect 5130 9215 5446 9216
rect 35850 9280 36166 9281
rect 35850 9216 35856 9280
rect 35920 9216 35936 9280
rect 36000 9216 36016 9280
rect 36080 9216 36096 9280
rect 36160 9216 36166 9280
rect 35850 9215 36166 9216
rect 66570 9280 66886 9281
rect 66570 9216 66576 9280
rect 66640 9216 66656 9280
rect 66720 9216 66736 9280
rect 66800 9216 66816 9280
rect 66880 9216 66886 9280
rect 66570 9215 66886 9216
rect 5790 8736 6106 8737
rect 5790 8672 5796 8736
rect 5860 8672 5876 8736
rect 5940 8672 5956 8736
rect 6020 8672 6036 8736
rect 6100 8672 6106 8736
rect 5790 8671 6106 8672
rect 36510 8736 36826 8737
rect 36510 8672 36516 8736
rect 36580 8672 36596 8736
rect 36660 8672 36676 8736
rect 36740 8672 36756 8736
rect 36820 8672 36826 8736
rect 36510 8671 36826 8672
rect 67230 8736 67546 8737
rect 67230 8672 67236 8736
rect 67300 8672 67316 8736
rect 67380 8672 67396 8736
rect 67460 8672 67476 8736
rect 67540 8672 67546 8736
rect 67230 8671 67546 8672
rect 5130 8192 5446 8193
rect 5130 8128 5136 8192
rect 5200 8128 5216 8192
rect 5280 8128 5296 8192
rect 5360 8128 5376 8192
rect 5440 8128 5446 8192
rect 5130 8127 5446 8128
rect 35850 8192 36166 8193
rect 35850 8128 35856 8192
rect 35920 8128 35936 8192
rect 36000 8128 36016 8192
rect 36080 8128 36096 8192
rect 36160 8128 36166 8192
rect 35850 8127 36166 8128
rect 66570 8192 66886 8193
rect 66570 8128 66576 8192
rect 66640 8128 66656 8192
rect 66720 8128 66736 8192
rect 66800 8128 66816 8192
rect 66880 8128 66886 8192
rect 66570 8127 66886 8128
rect 5790 7648 6106 7649
rect 5790 7584 5796 7648
rect 5860 7584 5876 7648
rect 5940 7584 5956 7648
rect 6020 7584 6036 7648
rect 6100 7584 6106 7648
rect 5790 7583 6106 7584
rect 36510 7648 36826 7649
rect 36510 7584 36516 7648
rect 36580 7584 36596 7648
rect 36660 7584 36676 7648
rect 36740 7584 36756 7648
rect 36820 7584 36826 7648
rect 36510 7583 36826 7584
rect 67230 7648 67546 7649
rect 67230 7584 67236 7648
rect 67300 7584 67316 7648
rect 67380 7584 67396 7648
rect 67460 7584 67476 7648
rect 67540 7584 67546 7648
rect 67230 7583 67546 7584
rect 5130 7104 5446 7105
rect 5130 7040 5136 7104
rect 5200 7040 5216 7104
rect 5280 7040 5296 7104
rect 5360 7040 5376 7104
rect 5440 7040 5446 7104
rect 5130 7039 5446 7040
rect 35850 7104 36166 7105
rect 35850 7040 35856 7104
rect 35920 7040 35936 7104
rect 36000 7040 36016 7104
rect 36080 7040 36096 7104
rect 36160 7040 36166 7104
rect 35850 7039 36166 7040
rect 66570 7104 66886 7105
rect 66570 7040 66576 7104
rect 66640 7040 66656 7104
rect 66720 7040 66736 7104
rect 66800 7040 66816 7104
rect 66880 7040 66886 7104
rect 66570 7039 66886 7040
rect 5790 6560 6106 6561
rect 5790 6496 5796 6560
rect 5860 6496 5876 6560
rect 5940 6496 5956 6560
rect 6020 6496 6036 6560
rect 6100 6496 6106 6560
rect 5790 6495 6106 6496
rect 36510 6560 36826 6561
rect 36510 6496 36516 6560
rect 36580 6496 36596 6560
rect 36660 6496 36676 6560
rect 36740 6496 36756 6560
rect 36820 6496 36826 6560
rect 36510 6495 36826 6496
rect 67230 6560 67546 6561
rect 67230 6496 67236 6560
rect 67300 6496 67316 6560
rect 67380 6496 67396 6560
rect 67460 6496 67476 6560
rect 67540 6496 67546 6560
rect 67230 6495 67546 6496
rect 5130 6016 5446 6017
rect 5130 5952 5136 6016
rect 5200 5952 5216 6016
rect 5280 5952 5296 6016
rect 5360 5952 5376 6016
rect 5440 5952 5446 6016
rect 5130 5951 5446 5952
rect 35850 6016 36166 6017
rect 35850 5952 35856 6016
rect 35920 5952 35936 6016
rect 36000 5952 36016 6016
rect 36080 5952 36096 6016
rect 36160 5952 36166 6016
rect 35850 5951 36166 5952
rect 66570 6016 66886 6017
rect 66570 5952 66576 6016
rect 66640 5952 66656 6016
rect 66720 5952 66736 6016
rect 66800 5952 66816 6016
rect 66880 5952 66886 6016
rect 66570 5951 66886 5952
rect 5790 5472 6106 5473
rect 5790 5408 5796 5472
rect 5860 5408 5876 5472
rect 5940 5408 5956 5472
rect 6020 5408 6036 5472
rect 6100 5408 6106 5472
rect 5790 5407 6106 5408
rect 36510 5472 36826 5473
rect 36510 5408 36516 5472
rect 36580 5408 36596 5472
rect 36660 5408 36676 5472
rect 36740 5408 36756 5472
rect 36820 5408 36826 5472
rect 36510 5407 36826 5408
rect 67230 5472 67546 5473
rect 67230 5408 67236 5472
rect 67300 5408 67316 5472
rect 67380 5408 67396 5472
rect 67460 5408 67476 5472
rect 67540 5408 67546 5472
rect 67230 5407 67546 5408
rect 5130 4928 5446 4929
rect 5130 4864 5136 4928
rect 5200 4864 5216 4928
rect 5280 4864 5296 4928
rect 5360 4864 5376 4928
rect 5440 4864 5446 4928
rect 5130 4863 5446 4864
rect 35850 4928 36166 4929
rect 35850 4864 35856 4928
rect 35920 4864 35936 4928
rect 36000 4864 36016 4928
rect 36080 4864 36096 4928
rect 36160 4864 36166 4928
rect 35850 4863 36166 4864
rect 66570 4928 66886 4929
rect 66570 4864 66576 4928
rect 66640 4864 66656 4928
rect 66720 4864 66736 4928
rect 66800 4864 66816 4928
rect 66880 4864 66886 4928
rect 66570 4863 66886 4864
rect 5790 4384 6106 4385
rect 5790 4320 5796 4384
rect 5860 4320 5876 4384
rect 5940 4320 5956 4384
rect 6020 4320 6036 4384
rect 6100 4320 6106 4384
rect 5790 4319 6106 4320
rect 36510 4384 36826 4385
rect 36510 4320 36516 4384
rect 36580 4320 36596 4384
rect 36660 4320 36676 4384
rect 36740 4320 36756 4384
rect 36820 4320 36826 4384
rect 36510 4319 36826 4320
rect 67230 4384 67546 4385
rect 67230 4320 67236 4384
rect 67300 4320 67316 4384
rect 67380 4320 67396 4384
rect 67460 4320 67476 4384
rect 67540 4320 67546 4384
rect 67230 4319 67546 4320
rect 5130 3840 5446 3841
rect 5130 3776 5136 3840
rect 5200 3776 5216 3840
rect 5280 3776 5296 3840
rect 5360 3776 5376 3840
rect 5440 3776 5446 3840
rect 5130 3775 5446 3776
rect 35850 3840 36166 3841
rect 35850 3776 35856 3840
rect 35920 3776 35936 3840
rect 36000 3776 36016 3840
rect 36080 3776 36096 3840
rect 36160 3776 36166 3840
rect 35850 3775 36166 3776
rect 66570 3840 66886 3841
rect 66570 3776 66576 3840
rect 66640 3776 66656 3840
rect 66720 3776 66736 3840
rect 66800 3776 66816 3840
rect 66880 3776 66886 3840
rect 66570 3775 66886 3776
rect 5790 3296 6106 3297
rect 5790 3232 5796 3296
rect 5860 3232 5876 3296
rect 5940 3232 5956 3296
rect 6020 3232 6036 3296
rect 6100 3232 6106 3296
rect 5790 3231 6106 3232
rect 36510 3296 36826 3297
rect 36510 3232 36516 3296
rect 36580 3232 36596 3296
rect 36660 3232 36676 3296
rect 36740 3232 36756 3296
rect 36820 3232 36826 3296
rect 36510 3231 36826 3232
rect 67230 3296 67546 3297
rect 67230 3232 67236 3296
rect 67300 3232 67316 3296
rect 67380 3232 67396 3296
rect 67460 3232 67476 3296
rect 67540 3232 67546 3296
rect 67230 3231 67546 3232
rect 5130 2752 5446 2753
rect 5130 2688 5136 2752
rect 5200 2688 5216 2752
rect 5280 2688 5296 2752
rect 5360 2688 5376 2752
rect 5440 2688 5446 2752
rect 5130 2687 5446 2688
rect 35850 2752 36166 2753
rect 35850 2688 35856 2752
rect 35920 2688 35936 2752
rect 36000 2688 36016 2752
rect 36080 2688 36096 2752
rect 36160 2688 36166 2752
rect 35850 2687 36166 2688
rect 66570 2752 66886 2753
rect 66570 2688 66576 2752
rect 66640 2688 66656 2752
rect 66720 2688 66736 2752
rect 66800 2688 66816 2752
rect 66880 2688 66886 2752
rect 66570 2687 66886 2688
rect 5790 2208 6106 2209
rect 5790 2144 5796 2208
rect 5860 2144 5876 2208
rect 5940 2144 5956 2208
rect 6020 2144 6036 2208
rect 6100 2144 6106 2208
rect 5790 2143 6106 2144
rect 36510 2208 36826 2209
rect 36510 2144 36516 2208
rect 36580 2144 36596 2208
rect 36660 2144 36676 2208
rect 36740 2144 36756 2208
rect 36820 2144 36826 2208
rect 36510 2143 36826 2144
rect 67230 2208 67546 2209
rect 67230 2144 67236 2208
rect 67300 2144 67316 2208
rect 67380 2144 67396 2208
rect 67460 2144 67476 2208
rect 67540 2144 67546 2208
rect 67230 2143 67546 2144
<< via3 >>
rect 5136 77820 5200 77824
rect 5136 77764 5140 77820
rect 5140 77764 5196 77820
rect 5196 77764 5200 77820
rect 5136 77760 5200 77764
rect 5216 77820 5280 77824
rect 5216 77764 5220 77820
rect 5220 77764 5276 77820
rect 5276 77764 5280 77820
rect 5216 77760 5280 77764
rect 5296 77820 5360 77824
rect 5296 77764 5300 77820
rect 5300 77764 5356 77820
rect 5356 77764 5360 77820
rect 5296 77760 5360 77764
rect 5376 77820 5440 77824
rect 5376 77764 5380 77820
rect 5380 77764 5436 77820
rect 5436 77764 5440 77820
rect 5376 77760 5440 77764
rect 35856 77820 35920 77824
rect 35856 77764 35860 77820
rect 35860 77764 35916 77820
rect 35916 77764 35920 77820
rect 35856 77760 35920 77764
rect 35936 77820 36000 77824
rect 35936 77764 35940 77820
rect 35940 77764 35996 77820
rect 35996 77764 36000 77820
rect 35936 77760 36000 77764
rect 36016 77820 36080 77824
rect 36016 77764 36020 77820
rect 36020 77764 36076 77820
rect 36076 77764 36080 77820
rect 36016 77760 36080 77764
rect 36096 77820 36160 77824
rect 36096 77764 36100 77820
rect 36100 77764 36156 77820
rect 36156 77764 36160 77820
rect 36096 77760 36160 77764
rect 66576 77820 66640 77824
rect 66576 77764 66580 77820
rect 66580 77764 66636 77820
rect 66636 77764 66640 77820
rect 66576 77760 66640 77764
rect 66656 77820 66720 77824
rect 66656 77764 66660 77820
rect 66660 77764 66716 77820
rect 66716 77764 66720 77820
rect 66656 77760 66720 77764
rect 66736 77820 66800 77824
rect 66736 77764 66740 77820
rect 66740 77764 66796 77820
rect 66796 77764 66800 77820
rect 66736 77760 66800 77764
rect 66816 77820 66880 77824
rect 66816 77764 66820 77820
rect 66820 77764 66876 77820
rect 66876 77764 66880 77820
rect 66816 77760 66880 77764
rect 5796 77276 5860 77280
rect 5796 77220 5800 77276
rect 5800 77220 5856 77276
rect 5856 77220 5860 77276
rect 5796 77216 5860 77220
rect 5876 77276 5940 77280
rect 5876 77220 5880 77276
rect 5880 77220 5936 77276
rect 5936 77220 5940 77276
rect 5876 77216 5940 77220
rect 5956 77276 6020 77280
rect 5956 77220 5960 77276
rect 5960 77220 6016 77276
rect 6016 77220 6020 77276
rect 5956 77216 6020 77220
rect 6036 77276 6100 77280
rect 6036 77220 6040 77276
rect 6040 77220 6096 77276
rect 6096 77220 6100 77276
rect 6036 77216 6100 77220
rect 36516 77276 36580 77280
rect 36516 77220 36520 77276
rect 36520 77220 36576 77276
rect 36576 77220 36580 77276
rect 36516 77216 36580 77220
rect 36596 77276 36660 77280
rect 36596 77220 36600 77276
rect 36600 77220 36656 77276
rect 36656 77220 36660 77276
rect 36596 77216 36660 77220
rect 36676 77276 36740 77280
rect 36676 77220 36680 77276
rect 36680 77220 36736 77276
rect 36736 77220 36740 77276
rect 36676 77216 36740 77220
rect 36756 77276 36820 77280
rect 36756 77220 36760 77276
rect 36760 77220 36816 77276
rect 36816 77220 36820 77276
rect 36756 77216 36820 77220
rect 67236 77276 67300 77280
rect 67236 77220 67240 77276
rect 67240 77220 67296 77276
rect 67296 77220 67300 77276
rect 67236 77216 67300 77220
rect 67316 77276 67380 77280
rect 67316 77220 67320 77276
rect 67320 77220 67376 77276
rect 67376 77220 67380 77276
rect 67316 77216 67380 77220
rect 67396 77276 67460 77280
rect 67396 77220 67400 77276
rect 67400 77220 67456 77276
rect 67456 77220 67460 77276
rect 67396 77216 67460 77220
rect 67476 77276 67540 77280
rect 67476 77220 67480 77276
rect 67480 77220 67536 77276
rect 67536 77220 67540 77276
rect 67476 77216 67540 77220
rect 5136 76732 5200 76736
rect 5136 76676 5140 76732
rect 5140 76676 5196 76732
rect 5196 76676 5200 76732
rect 5136 76672 5200 76676
rect 5216 76732 5280 76736
rect 5216 76676 5220 76732
rect 5220 76676 5276 76732
rect 5276 76676 5280 76732
rect 5216 76672 5280 76676
rect 5296 76732 5360 76736
rect 5296 76676 5300 76732
rect 5300 76676 5356 76732
rect 5356 76676 5360 76732
rect 5296 76672 5360 76676
rect 5376 76732 5440 76736
rect 5376 76676 5380 76732
rect 5380 76676 5436 76732
rect 5436 76676 5440 76732
rect 5376 76672 5440 76676
rect 35856 76732 35920 76736
rect 35856 76676 35860 76732
rect 35860 76676 35916 76732
rect 35916 76676 35920 76732
rect 35856 76672 35920 76676
rect 35936 76732 36000 76736
rect 35936 76676 35940 76732
rect 35940 76676 35996 76732
rect 35996 76676 36000 76732
rect 35936 76672 36000 76676
rect 36016 76732 36080 76736
rect 36016 76676 36020 76732
rect 36020 76676 36076 76732
rect 36076 76676 36080 76732
rect 36016 76672 36080 76676
rect 36096 76732 36160 76736
rect 36096 76676 36100 76732
rect 36100 76676 36156 76732
rect 36156 76676 36160 76732
rect 36096 76672 36160 76676
rect 66576 76732 66640 76736
rect 66576 76676 66580 76732
rect 66580 76676 66636 76732
rect 66636 76676 66640 76732
rect 66576 76672 66640 76676
rect 66656 76732 66720 76736
rect 66656 76676 66660 76732
rect 66660 76676 66716 76732
rect 66716 76676 66720 76732
rect 66656 76672 66720 76676
rect 66736 76732 66800 76736
rect 66736 76676 66740 76732
rect 66740 76676 66796 76732
rect 66796 76676 66800 76732
rect 66736 76672 66800 76676
rect 66816 76732 66880 76736
rect 66816 76676 66820 76732
rect 66820 76676 66876 76732
rect 66876 76676 66880 76732
rect 66816 76672 66880 76676
rect 5796 76188 5860 76192
rect 5796 76132 5800 76188
rect 5800 76132 5856 76188
rect 5856 76132 5860 76188
rect 5796 76128 5860 76132
rect 5876 76188 5940 76192
rect 5876 76132 5880 76188
rect 5880 76132 5936 76188
rect 5936 76132 5940 76188
rect 5876 76128 5940 76132
rect 5956 76188 6020 76192
rect 5956 76132 5960 76188
rect 5960 76132 6016 76188
rect 6016 76132 6020 76188
rect 5956 76128 6020 76132
rect 6036 76188 6100 76192
rect 6036 76132 6040 76188
rect 6040 76132 6096 76188
rect 6096 76132 6100 76188
rect 6036 76128 6100 76132
rect 36516 76188 36580 76192
rect 36516 76132 36520 76188
rect 36520 76132 36576 76188
rect 36576 76132 36580 76188
rect 36516 76128 36580 76132
rect 36596 76188 36660 76192
rect 36596 76132 36600 76188
rect 36600 76132 36656 76188
rect 36656 76132 36660 76188
rect 36596 76128 36660 76132
rect 36676 76188 36740 76192
rect 36676 76132 36680 76188
rect 36680 76132 36736 76188
rect 36736 76132 36740 76188
rect 36676 76128 36740 76132
rect 36756 76188 36820 76192
rect 36756 76132 36760 76188
rect 36760 76132 36816 76188
rect 36816 76132 36820 76188
rect 36756 76128 36820 76132
rect 67236 76188 67300 76192
rect 67236 76132 67240 76188
rect 67240 76132 67296 76188
rect 67296 76132 67300 76188
rect 67236 76128 67300 76132
rect 67316 76188 67380 76192
rect 67316 76132 67320 76188
rect 67320 76132 67376 76188
rect 67376 76132 67380 76188
rect 67316 76128 67380 76132
rect 67396 76188 67460 76192
rect 67396 76132 67400 76188
rect 67400 76132 67456 76188
rect 67456 76132 67460 76188
rect 67396 76128 67460 76132
rect 67476 76188 67540 76192
rect 67476 76132 67480 76188
rect 67480 76132 67536 76188
rect 67536 76132 67540 76188
rect 67476 76128 67540 76132
rect 5136 75644 5200 75648
rect 5136 75588 5140 75644
rect 5140 75588 5196 75644
rect 5196 75588 5200 75644
rect 5136 75584 5200 75588
rect 5216 75644 5280 75648
rect 5216 75588 5220 75644
rect 5220 75588 5276 75644
rect 5276 75588 5280 75644
rect 5216 75584 5280 75588
rect 5296 75644 5360 75648
rect 5296 75588 5300 75644
rect 5300 75588 5356 75644
rect 5356 75588 5360 75644
rect 5296 75584 5360 75588
rect 5376 75644 5440 75648
rect 5376 75588 5380 75644
rect 5380 75588 5436 75644
rect 5436 75588 5440 75644
rect 5376 75584 5440 75588
rect 35856 75644 35920 75648
rect 35856 75588 35860 75644
rect 35860 75588 35916 75644
rect 35916 75588 35920 75644
rect 35856 75584 35920 75588
rect 35936 75644 36000 75648
rect 35936 75588 35940 75644
rect 35940 75588 35996 75644
rect 35996 75588 36000 75644
rect 35936 75584 36000 75588
rect 36016 75644 36080 75648
rect 36016 75588 36020 75644
rect 36020 75588 36076 75644
rect 36076 75588 36080 75644
rect 36016 75584 36080 75588
rect 36096 75644 36160 75648
rect 36096 75588 36100 75644
rect 36100 75588 36156 75644
rect 36156 75588 36160 75644
rect 36096 75584 36160 75588
rect 66576 75644 66640 75648
rect 66576 75588 66580 75644
rect 66580 75588 66636 75644
rect 66636 75588 66640 75644
rect 66576 75584 66640 75588
rect 66656 75644 66720 75648
rect 66656 75588 66660 75644
rect 66660 75588 66716 75644
rect 66716 75588 66720 75644
rect 66656 75584 66720 75588
rect 66736 75644 66800 75648
rect 66736 75588 66740 75644
rect 66740 75588 66796 75644
rect 66796 75588 66800 75644
rect 66736 75584 66800 75588
rect 66816 75644 66880 75648
rect 66816 75588 66820 75644
rect 66820 75588 66876 75644
rect 66876 75588 66880 75644
rect 66816 75584 66880 75588
rect 5796 75100 5860 75104
rect 5796 75044 5800 75100
rect 5800 75044 5856 75100
rect 5856 75044 5860 75100
rect 5796 75040 5860 75044
rect 5876 75100 5940 75104
rect 5876 75044 5880 75100
rect 5880 75044 5936 75100
rect 5936 75044 5940 75100
rect 5876 75040 5940 75044
rect 5956 75100 6020 75104
rect 5956 75044 5960 75100
rect 5960 75044 6016 75100
rect 6016 75044 6020 75100
rect 5956 75040 6020 75044
rect 6036 75100 6100 75104
rect 6036 75044 6040 75100
rect 6040 75044 6096 75100
rect 6096 75044 6100 75100
rect 6036 75040 6100 75044
rect 36516 75100 36580 75104
rect 36516 75044 36520 75100
rect 36520 75044 36576 75100
rect 36576 75044 36580 75100
rect 36516 75040 36580 75044
rect 36596 75100 36660 75104
rect 36596 75044 36600 75100
rect 36600 75044 36656 75100
rect 36656 75044 36660 75100
rect 36596 75040 36660 75044
rect 36676 75100 36740 75104
rect 36676 75044 36680 75100
rect 36680 75044 36736 75100
rect 36736 75044 36740 75100
rect 36676 75040 36740 75044
rect 36756 75100 36820 75104
rect 36756 75044 36760 75100
rect 36760 75044 36816 75100
rect 36816 75044 36820 75100
rect 36756 75040 36820 75044
rect 67236 75100 67300 75104
rect 67236 75044 67240 75100
rect 67240 75044 67296 75100
rect 67296 75044 67300 75100
rect 67236 75040 67300 75044
rect 67316 75100 67380 75104
rect 67316 75044 67320 75100
rect 67320 75044 67376 75100
rect 67376 75044 67380 75100
rect 67316 75040 67380 75044
rect 67396 75100 67460 75104
rect 67396 75044 67400 75100
rect 67400 75044 67456 75100
rect 67456 75044 67460 75100
rect 67396 75040 67460 75044
rect 67476 75100 67540 75104
rect 67476 75044 67480 75100
rect 67480 75044 67536 75100
rect 67536 75044 67540 75100
rect 67476 75040 67540 75044
rect 5136 74556 5200 74560
rect 5136 74500 5140 74556
rect 5140 74500 5196 74556
rect 5196 74500 5200 74556
rect 5136 74496 5200 74500
rect 5216 74556 5280 74560
rect 5216 74500 5220 74556
rect 5220 74500 5276 74556
rect 5276 74500 5280 74556
rect 5216 74496 5280 74500
rect 5296 74556 5360 74560
rect 5296 74500 5300 74556
rect 5300 74500 5356 74556
rect 5356 74500 5360 74556
rect 5296 74496 5360 74500
rect 5376 74556 5440 74560
rect 5376 74500 5380 74556
rect 5380 74500 5436 74556
rect 5436 74500 5440 74556
rect 5376 74496 5440 74500
rect 35856 74556 35920 74560
rect 35856 74500 35860 74556
rect 35860 74500 35916 74556
rect 35916 74500 35920 74556
rect 35856 74496 35920 74500
rect 35936 74556 36000 74560
rect 35936 74500 35940 74556
rect 35940 74500 35996 74556
rect 35996 74500 36000 74556
rect 35936 74496 36000 74500
rect 36016 74556 36080 74560
rect 36016 74500 36020 74556
rect 36020 74500 36076 74556
rect 36076 74500 36080 74556
rect 36016 74496 36080 74500
rect 36096 74556 36160 74560
rect 36096 74500 36100 74556
rect 36100 74500 36156 74556
rect 36156 74500 36160 74556
rect 36096 74496 36160 74500
rect 66576 74556 66640 74560
rect 66576 74500 66580 74556
rect 66580 74500 66636 74556
rect 66636 74500 66640 74556
rect 66576 74496 66640 74500
rect 66656 74556 66720 74560
rect 66656 74500 66660 74556
rect 66660 74500 66716 74556
rect 66716 74500 66720 74556
rect 66656 74496 66720 74500
rect 66736 74556 66800 74560
rect 66736 74500 66740 74556
rect 66740 74500 66796 74556
rect 66796 74500 66800 74556
rect 66736 74496 66800 74500
rect 66816 74556 66880 74560
rect 66816 74500 66820 74556
rect 66820 74500 66876 74556
rect 66876 74500 66880 74556
rect 66816 74496 66880 74500
rect 5796 74012 5860 74016
rect 5796 73956 5800 74012
rect 5800 73956 5856 74012
rect 5856 73956 5860 74012
rect 5796 73952 5860 73956
rect 5876 74012 5940 74016
rect 5876 73956 5880 74012
rect 5880 73956 5936 74012
rect 5936 73956 5940 74012
rect 5876 73952 5940 73956
rect 5956 74012 6020 74016
rect 5956 73956 5960 74012
rect 5960 73956 6016 74012
rect 6016 73956 6020 74012
rect 5956 73952 6020 73956
rect 6036 74012 6100 74016
rect 6036 73956 6040 74012
rect 6040 73956 6096 74012
rect 6096 73956 6100 74012
rect 6036 73952 6100 73956
rect 36516 74012 36580 74016
rect 36516 73956 36520 74012
rect 36520 73956 36576 74012
rect 36576 73956 36580 74012
rect 36516 73952 36580 73956
rect 36596 74012 36660 74016
rect 36596 73956 36600 74012
rect 36600 73956 36656 74012
rect 36656 73956 36660 74012
rect 36596 73952 36660 73956
rect 36676 74012 36740 74016
rect 36676 73956 36680 74012
rect 36680 73956 36736 74012
rect 36736 73956 36740 74012
rect 36676 73952 36740 73956
rect 36756 74012 36820 74016
rect 36756 73956 36760 74012
rect 36760 73956 36816 74012
rect 36816 73956 36820 74012
rect 36756 73952 36820 73956
rect 67236 74012 67300 74016
rect 67236 73956 67240 74012
rect 67240 73956 67296 74012
rect 67296 73956 67300 74012
rect 67236 73952 67300 73956
rect 67316 74012 67380 74016
rect 67316 73956 67320 74012
rect 67320 73956 67376 74012
rect 67376 73956 67380 74012
rect 67316 73952 67380 73956
rect 67396 74012 67460 74016
rect 67396 73956 67400 74012
rect 67400 73956 67456 74012
rect 67456 73956 67460 74012
rect 67396 73952 67460 73956
rect 67476 74012 67540 74016
rect 67476 73956 67480 74012
rect 67480 73956 67536 74012
rect 67536 73956 67540 74012
rect 67476 73952 67540 73956
rect 5136 73468 5200 73472
rect 5136 73412 5140 73468
rect 5140 73412 5196 73468
rect 5196 73412 5200 73468
rect 5136 73408 5200 73412
rect 5216 73468 5280 73472
rect 5216 73412 5220 73468
rect 5220 73412 5276 73468
rect 5276 73412 5280 73468
rect 5216 73408 5280 73412
rect 5296 73468 5360 73472
rect 5296 73412 5300 73468
rect 5300 73412 5356 73468
rect 5356 73412 5360 73468
rect 5296 73408 5360 73412
rect 5376 73468 5440 73472
rect 5376 73412 5380 73468
rect 5380 73412 5436 73468
rect 5436 73412 5440 73468
rect 5376 73408 5440 73412
rect 35856 73468 35920 73472
rect 35856 73412 35860 73468
rect 35860 73412 35916 73468
rect 35916 73412 35920 73468
rect 35856 73408 35920 73412
rect 35936 73468 36000 73472
rect 35936 73412 35940 73468
rect 35940 73412 35996 73468
rect 35996 73412 36000 73468
rect 35936 73408 36000 73412
rect 36016 73468 36080 73472
rect 36016 73412 36020 73468
rect 36020 73412 36076 73468
rect 36076 73412 36080 73468
rect 36016 73408 36080 73412
rect 36096 73468 36160 73472
rect 36096 73412 36100 73468
rect 36100 73412 36156 73468
rect 36156 73412 36160 73468
rect 36096 73408 36160 73412
rect 66576 73468 66640 73472
rect 66576 73412 66580 73468
rect 66580 73412 66636 73468
rect 66636 73412 66640 73468
rect 66576 73408 66640 73412
rect 66656 73468 66720 73472
rect 66656 73412 66660 73468
rect 66660 73412 66716 73468
rect 66716 73412 66720 73468
rect 66656 73408 66720 73412
rect 66736 73468 66800 73472
rect 66736 73412 66740 73468
rect 66740 73412 66796 73468
rect 66796 73412 66800 73468
rect 66736 73408 66800 73412
rect 66816 73468 66880 73472
rect 66816 73412 66820 73468
rect 66820 73412 66876 73468
rect 66876 73412 66880 73468
rect 66816 73408 66880 73412
rect 5796 72924 5860 72928
rect 5796 72868 5800 72924
rect 5800 72868 5856 72924
rect 5856 72868 5860 72924
rect 5796 72864 5860 72868
rect 5876 72924 5940 72928
rect 5876 72868 5880 72924
rect 5880 72868 5936 72924
rect 5936 72868 5940 72924
rect 5876 72864 5940 72868
rect 5956 72924 6020 72928
rect 5956 72868 5960 72924
rect 5960 72868 6016 72924
rect 6016 72868 6020 72924
rect 5956 72864 6020 72868
rect 6036 72924 6100 72928
rect 6036 72868 6040 72924
rect 6040 72868 6096 72924
rect 6096 72868 6100 72924
rect 6036 72864 6100 72868
rect 36516 72924 36580 72928
rect 36516 72868 36520 72924
rect 36520 72868 36576 72924
rect 36576 72868 36580 72924
rect 36516 72864 36580 72868
rect 36596 72924 36660 72928
rect 36596 72868 36600 72924
rect 36600 72868 36656 72924
rect 36656 72868 36660 72924
rect 36596 72864 36660 72868
rect 36676 72924 36740 72928
rect 36676 72868 36680 72924
rect 36680 72868 36736 72924
rect 36736 72868 36740 72924
rect 36676 72864 36740 72868
rect 36756 72924 36820 72928
rect 36756 72868 36760 72924
rect 36760 72868 36816 72924
rect 36816 72868 36820 72924
rect 36756 72864 36820 72868
rect 67236 72924 67300 72928
rect 67236 72868 67240 72924
rect 67240 72868 67296 72924
rect 67296 72868 67300 72924
rect 67236 72864 67300 72868
rect 67316 72924 67380 72928
rect 67316 72868 67320 72924
rect 67320 72868 67376 72924
rect 67376 72868 67380 72924
rect 67316 72864 67380 72868
rect 67396 72924 67460 72928
rect 67396 72868 67400 72924
rect 67400 72868 67456 72924
rect 67456 72868 67460 72924
rect 67396 72864 67460 72868
rect 67476 72924 67540 72928
rect 67476 72868 67480 72924
rect 67480 72868 67536 72924
rect 67536 72868 67540 72924
rect 67476 72864 67540 72868
rect 5136 72380 5200 72384
rect 5136 72324 5140 72380
rect 5140 72324 5196 72380
rect 5196 72324 5200 72380
rect 5136 72320 5200 72324
rect 5216 72380 5280 72384
rect 5216 72324 5220 72380
rect 5220 72324 5276 72380
rect 5276 72324 5280 72380
rect 5216 72320 5280 72324
rect 5296 72380 5360 72384
rect 5296 72324 5300 72380
rect 5300 72324 5356 72380
rect 5356 72324 5360 72380
rect 5296 72320 5360 72324
rect 5376 72380 5440 72384
rect 5376 72324 5380 72380
rect 5380 72324 5436 72380
rect 5436 72324 5440 72380
rect 5376 72320 5440 72324
rect 35856 72380 35920 72384
rect 35856 72324 35860 72380
rect 35860 72324 35916 72380
rect 35916 72324 35920 72380
rect 35856 72320 35920 72324
rect 35936 72380 36000 72384
rect 35936 72324 35940 72380
rect 35940 72324 35996 72380
rect 35996 72324 36000 72380
rect 35936 72320 36000 72324
rect 36016 72380 36080 72384
rect 36016 72324 36020 72380
rect 36020 72324 36076 72380
rect 36076 72324 36080 72380
rect 36016 72320 36080 72324
rect 36096 72380 36160 72384
rect 36096 72324 36100 72380
rect 36100 72324 36156 72380
rect 36156 72324 36160 72380
rect 36096 72320 36160 72324
rect 66576 72380 66640 72384
rect 66576 72324 66580 72380
rect 66580 72324 66636 72380
rect 66636 72324 66640 72380
rect 66576 72320 66640 72324
rect 66656 72380 66720 72384
rect 66656 72324 66660 72380
rect 66660 72324 66716 72380
rect 66716 72324 66720 72380
rect 66656 72320 66720 72324
rect 66736 72380 66800 72384
rect 66736 72324 66740 72380
rect 66740 72324 66796 72380
rect 66796 72324 66800 72380
rect 66736 72320 66800 72324
rect 66816 72380 66880 72384
rect 66816 72324 66820 72380
rect 66820 72324 66876 72380
rect 66876 72324 66880 72380
rect 66816 72320 66880 72324
rect 5796 71836 5860 71840
rect 5796 71780 5800 71836
rect 5800 71780 5856 71836
rect 5856 71780 5860 71836
rect 5796 71776 5860 71780
rect 5876 71836 5940 71840
rect 5876 71780 5880 71836
rect 5880 71780 5936 71836
rect 5936 71780 5940 71836
rect 5876 71776 5940 71780
rect 5956 71836 6020 71840
rect 5956 71780 5960 71836
rect 5960 71780 6016 71836
rect 6016 71780 6020 71836
rect 5956 71776 6020 71780
rect 6036 71836 6100 71840
rect 6036 71780 6040 71836
rect 6040 71780 6096 71836
rect 6096 71780 6100 71836
rect 6036 71776 6100 71780
rect 36516 71836 36580 71840
rect 36516 71780 36520 71836
rect 36520 71780 36576 71836
rect 36576 71780 36580 71836
rect 36516 71776 36580 71780
rect 36596 71836 36660 71840
rect 36596 71780 36600 71836
rect 36600 71780 36656 71836
rect 36656 71780 36660 71836
rect 36596 71776 36660 71780
rect 36676 71836 36740 71840
rect 36676 71780 36680 71836
rect 36680 71780 36736 71836
rect 36736 71780 36740 71836
rect 36676 71776 36740 71780
rect 36756 71836 36820 71840
rect 36756 71780 36760 71836
rect 36760 71780 36816 71836
rect 36816 71780 36820 71836
rect 36756 71776 36820 71780
rect 67236 71836 67300 71840
rect 67236 71780 67240 71836
rect 67240 71780 67296 71836
rect 67296 71780 67300 71836
rect 67236 71776 67300 71780
rect 67316 71836 67380 71840
rect 67316 71780 67320 71836
rect 67320 71780 67376 71836
rect 67376 71780 67380 71836
rect 67316 71776 67380 71780
rect 67396 71836 67460 71840
rect 67396 71780 67400 71836
rect 67400 71780 67456 71836
rect 67456 71780 67460 71836
rect 67396 71776 67460 71780
rect 67476 71836 67540 71840
rect 67476 71780 67480 71836
rect 67480 71780 67536 71836
rect 67536 71780 67540 71836
rect 67476 71776 67540 71780
rect 5136 71292 5200 71296
rect 5136 71236 5140 71292
rect 5140 71236 5196 71292
rect 5196 71236 5200 71292
rect 5136 71232 5200 71236
rect 5216 71292 5280 71296
rect 5216 71236 5220 71292
rect 5220 71236 5276 71292
rect 5276 71236 5280 71292
rect 5216 71232 5280 71236
rect 5296 71292 5360 71296
rect 5296 71236 5300 71292
rect 5300 71236 5356 71292
rect 5356 71236 5360 71292
rect 5296 71232 5360 71236
rect 5376 71292 5440 71296
rect 5376 71236 5380 71292
rect 5380 71236 5436 71292
rect 5436 71236 5440 71292
rect 5376 71232 5440 71236
rect 35856 71292 35920 71296
rect 35856 71236 35860 71292
rect 35860 71236 35916 71292
rect 35916 71236 35920 71292
rect 35856 71232 35920 71236
rect 35936 71292 36000 71296
rect 35936 71236 35940 71292
rect 35940 71236 35996 71292
rect 35996 71236 36000 71292
rect 35936 71232 36000 71236
rect 36016 71292 36080 71296
rect 36016 71236 36020 71292
rect 36020 71236 36076 71292
rect 36076 71236 36080 71292
rect 36016 71232 36080 71236
rect 36096 71292 36160 71296
rect 36096 71236 36100 71292
rect 36100 71236 36156 71292
rect 36156 71236 36160 71292
rect 36096 71232 36160 71236
rect 66576 71292 66640 71296
rect 66576 71236 66580 71292
rect 66580 71236 66636 71292
rect 66636 71236 66640 71292
rect 66576 71232 66640 71236
rect 66656 71292 66720 71296
rect 66656 71236 66660 71292
rect 66660 71236 66716 71292
rect 66716 71236 66720 71292
rect 66656 71232 66720 71236
rect 66736 71292 66800 71296
rect 66736 71236 66740 71292
rect 66740 71236 66796 71292
rect 66796 71236 66800 71292
rect 66736 71232 66800 71236
rect 66816 71292 66880 71296
rect 66816 71236 66820 71292
rect 66820 71236 66876 71292
rect 66876 71236 66880 71292
rect 66816 71232 66880 71236
rect 5796 70748 5860 70752
rect 5796 70692 5800 70748
rect 5800 70692 5856 70748
rect 5856 70692 5860 70748
rect 5796 70688 5860 70692
rect 5876 70748 5940 70752
rect 5876 70692 5880 70748
rect 5880 70692 5936 70748
rect 5936 70692 5940 70748
rect 5876 70688 5940 70692
rect 5956 70748 6020 70752
rect 5956 70692 5960 70748
rect 5960 70692 6016 70748
rect 6016 70692 6020 70748
rect 5956 70688 6020 70692
rect 6036 70748 6100 70752
rect 6036 70692 6040 70748
rect 6040 70692 6096 70748
rect 6096 70692 6100 70748
rect 6036 70688 6100 70692
rect 36516 70748 36580 70752
rect 36516 70692 36520 70748
rect 36520 70692 36576 70748
rect 36576 70692 36580 70748
rect 36516 70688 36580 70692
rect 36596 70748 36660 70752
rect 36596 70692 36600 70748
rect 36600 70692 36656 70748
rect 36656 70692 36660 70748
rect 36596 70688 36660 70692
rect 36676 70748 36740 70752
rect 36676 70692 36680 70748
rect 36680 70692 36736 70748
rect 36736 70692 36740 70748
rect 36676 70688 36740 70692
rect 36756 70748 36820 70752
rect 36756 70692 36760 70748
rect 36760 70692 36816 70748
rect 36816 70692 36820 70748
rect 36756 70688 36820 70692
rect 67236 70748 67300 70752
rect 67236 70692 67240 70748
rect 67240 70692 67296 70748
rect 67296 70692 67300 70748
rect 67236 70688 67300 70692
rect 67316 70748 67380 70752
rect 67316 70692 67320 70748
rect 67320 70692 67376 70748
rect 67376 70692 67380 70748
rect 67316 70688 67380 70692
rect 67396 70748 67460 70752
rect 67396 70692 67400 70748
rect 67400 70692 67456 70748
rect 67456 70692 67460 70748
rect 67396 70688 67460 70692
rect 67476 70748 67540 70752
rect 67476 70692 67480 70748
rect 67480 70692 67536 70748
rect 67536 70692 67540 70748
rect 67476 70688 67540 70692
rect 5136 70204 5200 70208
rect 5136 70148 5140 70204
rect 5140 70148 5196 70204
rect 5196 70148 5200 70204
rect 5136 70144 5200 70148
rect 5216 70204 5280 70208
rect 5216 70148 5220 70204
rect 5220 70148 5276 70204
rect 5276 70148 5280 70204
rect 5216 70144 5280 70148
rect 5296 70204 5360 70208
rect 5296 70148 5300 70204
rect 5300 70148 5356 70204
rect 5356 70148 5360 70204
rect 5296 70144 5360 70148
rect 5376 70204 5440 70208
rect 5376 70148 5380 70204
rect 5380 70148 5436 70204
rect 5436 70148 5440 70204
rect 5376 70144 5440 70148
rect 35856 70204 35920 70208
rect 35856 70148 35860 70204
rect 35860 70148 35916 70204
rect 35916 70148 35920 70204
rect 35856 70144 35920 70148
rect 35936 70204 36000 70208
rect 35936 70148 35940 70204
rect 35940 70148 35996 70204
rect 35996 70148 36000 70204
rect 35936 70144 36000 70148
rect 36016 70204 36080 70208
rect 36016 70148 36020 70204
rect 36020 70148 36076 70204
rect 36076 70148 36080 70204
rect 36016 70144 36080 70148
rect 36096 70204 36160 70208
rect 36096 70148 36100 70204
rect 36100 70148 36156 70204
rect 36156 70148 36160 70204
rect 36096 70144 36160 70148
rect 66576 70204 66640 70208
rect 66576 70148 66580 70204
rect 66580 70148 66636 70204
rect 66636 70148 66640 70204
rect 66576 70144 66640 70148
rect 66656 70204 66720 70208
rect 66656 70148 66660 70204
rect 66660 70148 66716 70204
rect 66716 70148 66720 70204
rect 66656 70144 66720 70148
rect 66736 70204 66800 70208
rect 66736 70148 66740 70204
rect 66740 70148 66796 70204
rect 66796 70148 66800 70204
rect 66736 70144 66800 70148
rect 66816 70204 66880 70208
rect 66816 70148 66820 70204
rect 66820 70148 66876 70204
rect 66876 70148 66880 70204
rect 66816 70144 66880 70148
rect 5796 69660 5860 69664
rect 5796 69604 5800 69660
rect 5800 69604 5856 69660
rect 5856 69604 5860 69660
rect 5796 69600 5860 69604
rect 5876 69660 5940 69664
rect 5876 69604 5880 69660
rect 5880 69604 5936 69660
rect 5936 69604 5940 69660
rect 5876 69600 5940 69604
rect 5956 69660 6020 69664
rect 5956 69604 5960 69660
rect 5960 69604 6016 69660
rect 6016 69604 6020 69660
rect 5956 69600 6020 69604
rect 6036 69660 6100 69664
rect 6036 69604 6040 69660
rect 6040 69604 6096 69660
rect 6096 69604 6100 69660
rect 6036 69600 6100 69604
rect 36516 69660 36580 69664
rect 36516 69604 36520 69660
rect 36520 69604 36576 69660
rect 36576 69604 36580 69660
rect 36516 69600 36580 69604
rect 36596 69660 36660 69664
rect 36596 69604 36600 69660
rect 36600 69604 36656 69660
rect 36656 69604 36660 69660
rect 36596 69600 36660 69604
rect 36676 69660 36740 69664
rect 36676 69604 36680 69660
rect 36680 69604 36736 69660
rect 36736 69604 36740 69660
rect 36676 69600 36740 69604
rect 36756 69660 36820 69664
rect 36756 69604 36760 69660
rect 36760 69604 36816 69660
rect 36816 69604 36820 69660
rect 36756 69600 36820 69604
rect 67236 69660 67300 69664
rect 67236 69604 67240 69660
rect 67240 69604 67296 69660
rect 67296 69604 67300 69660
rect 67236 69600 67300 69604
rect 67316 69660 67380 69664
rect 67316 69604 67320 69660
rect 67320 69604 67376 69660
rect 67376 69604 67380 69660
rect 67316 69600 67380 69604
rect 67396 69660 67460 69664
rect 67396 69604 67400 69660
rect 67400 69604 67456 69660
rect 67456 69604 67460 69660
rect 67396 69600 67460 69604
rect 67476 69660 67540 69664
rect 67476 69604 67480 69660
rect 67480 69604 67536 69660
rect 67536 69604 67540 69660
rect 67476 69600 67540 69604
rect 5136 69116 5200 69120
rect 5136 69060 5140 69116
rect 5140 69060 5196 69116
rect 5196 69060 5200 69116
rect 5136 69056 5200 69060
rect 5216 69116 5280 69120
rect 5216 69060 5220 69116
rect 5220 69060 5276 69116
rect 5276 69060 5280 69116
rect 5216 69056 5280 69060
rect 5296 69116 5360 69120
rect 5296 69060 5300 69116
rect 5300 69060 5356 69116
rect 5356 69060 5360 69116
rect 5296 69056 5360 69060
rect 5376 69116 5440 69120
rect 5376 69060 5380 69116
rect 5380 69060 5436 69116
rect 5436 69060 5440 69116
rect 5376 69056 5440 69060
rect 35856 69116 35920 69120
rect 35856 69060 35860 69116
rect 35860 69060 35916 69116
rect 35916 69060 35920 69116
rect 35856 69056 35920 69060
rect 35936 69116 36000 69120
rect 35936 69060 35940 69116
rect 35940 69060 35996 69116
rect 35996 69060 36000 69116
rect 35936 69056 36000 69060
rect 36016 69116 36080 69120
rect 36016 69060 36020 69116
rect 36020 69060 36076 69116
rect 36076 69060 36080 69116
rect 36016 69056 36080 69060
rect 36096 69116 36160 69120
rect 36096 69060 36100 69116
rect 36100 69060 36156 69116
rect 36156 69060 36160 69116
rect 36096 69056 36160 69060
rect 66576 69116 66640 69120
rect 66576 69060 66580 69116
rect 66580 69060 66636 69116
rect 66636 69060 66640 69116
rect 66576 69056 66640 69060
rect 66656 69116 66720 69120
rect 66656 69060 66660 69116
rect 66660 69060 66716 69116
rect 66716 69060 66720 69116
rect 66656 69056 66720 69060
rect 66736 69116 66800 69120
rect 66736 69060 66740 69116
rect 66740 69060 66796 69116
rect 66796 69060 66800 69116
rect 66736 69056 66800 69060
rect 66816 69116 66880 69120
rect 66816 69060 66820 69116
rect 66820 69060 66876 69116
rect 66876 69060 66880 69116
rect 66816 69056 66880 69060
rect 5796 68572 5860 68576
rect 5796 68516 5800 68572
rect 5800 68516 5856 68572
rect 5856 68516 5860 68572
rect 5796 68512 5860 68516
rect 5876 68572 5940 68576
rect 5876 68516 5880 68572
rect 5880 68516 5936 68572
rect 5936 68516 5940 68572
rect 5876 68512 5940 68516
rect 5956 68572 6020 68576
rect 5956 68516 5960 68572
rect 5960 68516 6016 68572
rect 6016 68516 6020 68572
rect 5956 68512 6020 68516
rect 6036 68572 6100 68576
rect 6036 68516 6040 68572
rect 6040 68516 6096 68572
rect 6096 68516 6100 68572
rect 6036 68512 6100 68516
rect 36516 68572 36580 68576
rect 36516 68516 36520 68572
rect 36520 68516 36576 68572
rect 36576 68516 36580 68572
rect 36516 68512 36580 68516
rect 36596 68572 36660 68576
rect 36596 68516 36600 68572
rect 36600 68516 36656 68572
rect 36656 68516 36660 68572
rect 36596 68512 36660 68516
rect 36676 68572 36740 68576
rect 36676 68516 36680 68572
rect 36680 68516 36736 68572
rect 36736 68516 36740 68572
rect 36676 68512 36740 68516
rect 36756 68572 36820 68576
rect 36756 68516 36760 68572
rect 36760 68516 36816 68572
rect 36816 68516 36820 68572
rect 36756 68512 36820 68516
rect 67236 68572 67300 68576
rect 67236 68516 67240 68572
rect 67240 68516 67296 68572
rect 67296 68516 67300 68572
rect 67236 68512 67300 68516
rect 67316 68572 67380 68576
rect 67316 68516 67320 68572
rect 67320 68516 67376 68572
rect 67376 68516 67380 68572
rect 67316 68512 67380 68516
rect 67396 68572 67460 68576
rect 67396 68516 67400 68572
rect 67400 68516 67456 68572
rect 67456 68516 67460 68572
rect 67396 68512 67460 68516
rect 67476 68572 67540 68576
rect 67476 68516 67480 68572
rect 67480 68516 67536 68572
rect 67536 68516 67540 68572
rect 67476 68512 67540 68516
rect 5136 68028 5200 68032
rect 5136 67972 5140 68028
rect 5140 67972 5196 68028
rect 5196 67972 5200 68028
rect 5136 67968 5200 67972
rect 5216 68028 5280 68032
rect 5216 67972 5220 68028
rect 5220 67972 5276 68028
rect 5276 67972 5280 68028
rect 5216 67968 5280 67972
rect 5296 68028 5360 68032
rect 5296 67972 5300 68028
rect 5300 67972 5356 68028
rect 5356 67972 5360 68028
rect 5296 67968 5360 67972
rect 5376 68028 5440 68032
rect 5376 67972 5380 68028
rect 5380 67972 5436 68028
rect 5436 67972 5440 68028
rect 5376 67968 5440 67972
rect 35856 68028 35920 68032
rect 35856 67972 35860 68028
rect 35860 67972 35916 68028
rect 35916 67972 35920 68028
rect 35856 67968 35920 67972
rect 35936 68028 36000 68032
rect 35936 67972 35940 68028
rect 35940 67972 35996 68028
rect 35996 67972 36000 68028
rect 35936 67968 36000 67972
rect 36016 68028 36080 68032
rect 36016 67972 36020 68028
rect 36020 67972 36076 68028
rect 36076 67972 36080 68028
rect 36016 67968 36080 67972
rect 36096 68028 36160 68032
rect 36096 67972 36100 68028
rect 36100 67972 36156 68028
rect 36156 67972 36160 68028
rect 36096 67968 36160 67972
rect 66576 68028 66640 68032
rect 66576 67972 66580 68028
rect 66580 67972 66636 68028
rect 66636 67972 66640 68028
rect 66576 67968 66640 67972
rect 66656 68028 66720 68032
rect 66656 67972 66660 68028
rect 66660 67972 66716 68028
rect 66716 67972 66720 68028
rect 66656 67968 66720 67972
rect 66736 68028 66800 68032
rect 66736 67972 66740 68028
rect 66740 67972 66796 68028
rect 66796 67972 66800 68028
rect 66736 67968 66800 67972
rect 66816 68028 66880 68032
rect 66816 67972 66820 68028
rect 66820 67972 66876 68028
rect 66876 67972 66880 68028
rect 66816 67968 66880 67972
rect 5796 67484 5860 67488
rect 5796 67428 5800 67484
rect 5800 67428 5856 67484
rect 5856 67428 5860 67484
rect 5796 67424 5860 67428
rect 5876 67484 5940 67488
rect 5876 67428 5880 67484
rect 5880 67428 5936 67484
rect 5936 67428 5940 67484
rect 5876 67424 5940 67428
rect 5956 67484 6020 67488
rect 5956 67428 5960 67484
rect 5960 67428 6016 67484
rect 6016 67428 6020 67484
rect 5956 67424 6020 67428
rect 6036 67484 6100 67488
rect 6036 67428 6040 67484
rect 6040 67428 6096 67484
rect 6096 67428 6100 67484
rect 6036 67424 6100 67428
rect 36516 67484 36580 67488
rect 36516 67428 36520 67484
rect 36520 67428 36576 67484
rect 36576 67428 36580 67484
rect 36516 67424 36580 67428
rect 36596 67484 36660 67488
rect 36596 67428 36600 67484
rect 36600 67428 36656 67484
rect 36656 67428 36660 67484
rect 36596 67424 36660 67428
rect 36676 67484 36740 67488
rect 36676 67428 36680 67484
rect 36680 67428 36736 67484
rect 36736 67428 36740 67484
rect 36676 67424 36740 67428
rect 36756 67484 36820 67488
rect 36756 67428 36760 67484
rect 36760 67428 36816 67484
rect 36816 67428 36820 67484
rect 36756 67424 36820 67428
rect 67236 67484 67300 67488
rect 67236 67428 67240 67484
rect 67240 67428 67296 67484
rect 67296 67428 67300 67484
rect 67236 67424 67300 67428
rect 67316 67484 67380 67488
rect 67316 67428 67320 67484
rect 67320 67428 67376 67484
rect 67376 67428 67380 67484
rect 67316 67424 67380 67428
rect 67396 67484 67460 67488
rect 67396 67428 67400 67484
rect 67400 67428 67456 67484
rect 67456 67428 67460 67484
rect 67396 67424 67460 67428
rect 67476 67484 67540 67488
rect 67476 67428 67480 67484
rect 67480 67428 67536 67484
rect 67536 67428 67540 67484
rect 67476 67424 67540 67428
rect 5136 66940 5200 66944
rect 5136 66884 5140 66940
rect 5140 66884 5196 66940
rect 5196 66884 5200 66940
rect 5136 66880 5200 66884
rect 5216 66940 5280 66944
rect 5216 66884 5220 66940
rect 5220 66884 5276 66940
rect 5276 66884 5280 66940
rect 5216 66880 5280 66884
rect 5296 66940 5360 66944
rect 5296 66884 5300 66940
rect 5300 66884 5356 66940
rect 5356 66884 5360 66940
rect 5296 66880 5360 66884
rect 5376 66940 5440 66944
rect 5376 66884 5380 66940
rect 5380 66884 5436 66940
rect 5436 66884 5440 66940
rect 5376 66880 5440 66884
rect 35856 66940 35920 66944
rect 35856 66884 35860 66940
rect 35860 66884 35916 66940
rect 35916 66884 35920 66940
rect 35856 66880 35920 66884
rect 35936 66940 36000 66944
rect 35936 66884 35940 66940
rect 35940 66884 35996 66940
rect 35996 66884 36000 66940
rect 35936 66880 36000 66884
rect 36016 66940 36080 66944
rect 36016 66884 36020 66940
rect 36020 66884 36076 66940
rect 36076 66884 36080 66940
rect 36016 66880 36080 66884
rect 36096 66940 36160 66944
rect 36096 66884 36100 66940
rect 36100 66884 36156 66940
rect 36156 66884 36160 66940
rect 36096 66880 36160 66884
rect 66576 66940 66640 66944
rect 66576 66884 66580 66940
rect 66580 66884 66636 66940
rect 66636 66884 66640 66940
rect 66576 66880 66640 66884
rect 66656 66940 66720 66944
rect 66656 66884 66660 66940
rect 66660 66884 66716 66940
rect 66716 66884 66720 66940
rect 66656 66880 66720 66884
rect 66736 66940 66800 66944
rect 66736 66884 66740 66940
rect 66740 66884 66796 66940
rect 66796 66884 66800 66940
rect 66736 66880 66800 66884
rect 66816 66940 66880 66944
rect 66816 66884 66820 66940
rect 66820 66884 66876 66940
rect 66876 66884 66880 66940
rect 66816 66880 66880 66884
rect 5796 66396 5860 66400
rect 5796 66340 5800 66396
rect 5800 66340 5856 66396
rect 5856 66340 5860 66396
rect 5796 66336 5860 66340
rect 5876 66396 5940 66400
rect 5876 66340 5880 66396
rect 5880 66340 5936 66396
rect 5936 66340 5940 66396
rect 5876 66336 5940 66340
rect 5956 66396 6020 66400
rect 5956 66340 5960 66396
rect 5960 66340 6016 66396
rect 6016 66340 6020 66396
rect 5956 66336 6020 66340
rect 6036 66396 6100 66400
rect 6036 66340 6040 66396
rect 6040 66340 6096 66396
rect 6096 66340 6100 66396
rect 6036 66336 6100 66340
rect 36516 66396 36580 66400
rect 36516 66340 36520 66396
rect 36520 66340 36576 66396
rect 36576 66340 36580 66396
rect 36516 66336 36580 66340
rect 36596 66396 36660 66400
rect 36596 66340 36600 66396
rect 36600 66340 36656 66396
rect 36656 66340 36660 66396
rect 36596 66336 36660 66340
rect 36676 66396 36740 66400
rect 36676 66340 36680 66396
rect 36680 66340 36736 66396
rect 36736 66340 36740 66396
rect 36676 66336 36740 66340
rect 36756 66396 36820 66400
rect 36756 66340 36760 66396
rect 36760 66340 36816 66396
rect 36816 66340 36820 66396
rect 36756 66336 36820 66340
rect 67236 66396 67300 66400
rect 67236 66340 67240 66396
rect 67240 66340 67296 66396
rect 67296 66340 67300 66396
rect 67236 66336 67300 66340
rect 67316 66396 67380 66400
rect 67316 66340 67320 66396
rect 67320 66340 67376 66396
rect 67376 66340 67380 66396
rect 67316 66336 67380 66340
rect 67396 66396 67460 66400
rect 67396 66340 67400 66396
rect 67400 66340 67456 66396
rect 67456 66340 67460 66396
rect 67396 66336 67460 66340
rect 67476 66396 67540 66400
rect 67476 66340 67480 66396
rect 67480 66340 67536 66396
rect 67536 66340 67540 66396
rect 67476 66336 67540 66340
rect 5136 65852 5200 65856
rect 5136 65796 5140 65852
rect 5140 65796 5196 65852
rect 5196 65796 5200 65852
rect 5136 65792 5200 65796
rect 5216 65852 5280 65856
rect 5216 65796 5220 65852
rect 5220 65796 5276 65852
rect 5276 65796 5280 65852
rect 5216 65792 5280 65796
rect 5296 65852 5360 65856
rect 5296 65796 5300 65852
rect 5300 65796 5356 65852
rect 5356 65796 5360 65852
rect 5296 65792 5360 65796
rect 5376 65852 5440 65856
rect 5376 65796 5380 65852
rect 5380 65796 5436 65852
rect 5436 65796 5440 65852
rect 5376 65792 5440 65796
rect 35856 65852 35920 65856
rect 35856 65796 35860 65852
rect 35860 65796 35916 65852
rect 35916 65796 35920 65852
rect 35856 65792 35920 65796
rect 35936 65852 36000 65856
rect 35936 65796 35940 65852
rect 35940 65796 35996 65852
rect 35996 65796 36000 65852
rect 35936 65792 36000 65796
rect 36016 65852 36080 65856
rect 36016 65796 36020 65852
rect 36020 65796 36076 65852
rect 36076 65796 36080 65852
rect 36016 65792 36080 65796
rect 36096 65852 36160 65856
rect 36096 65796 36100 65852
rect 36100 65796 36156 65852
rect 36156 65796 36160 65852
rect 36096 65792 36160 65796
rect 66576 65852 66640 65856
rect 66576 65796 66580 65852
rect 66580 65796 66636 65852
rect 66636 65796 66640 65852
rect 66576 65792 66640 65796
rect 66656 65852 66720 65856
rect 66656 65796 66660 65852
rect 66660 65796 66716 65852
rect 66716 65796 66720 65852
rect 66656 65792 66720 65796
rect 66736 65852 66800 65856
rect 66736 65796 66740 65852
rect 66740 65796 66796 65852
rect 66796 65796 66800 65852
rect 66736 65792 66800 65796
rect 66816 65852 66880 65856
rect 66816 65796 66820 65852
rect 66820 65796 66876 65852
rect 66876 65796 66880 65852
rect 66816 65792 66880 65796
rect 5796 65308 5860 65312
rect 5796 65252 5800 65308
rect 5800 65252 5856 65308
rect 5856 65252 5860 65308
rect 5796 65248 5860 65252
rect 5876 65308 5940 65312
rect 5876 65252 5880 65308
rect 5880 65252 5936 65308
rect 5936 65252 5940 65308
rect 5876 65248 5940 65252
rect 5956 65308 6020 65312
rect 5956 65252 5960 65308
rect 5960 65252 6016 65308
rect 6016 65252 6020 65308
rect 5956 65248 6020 65252
rect 6036 65308 6100 65312
rect 6036 65252 6040 65308
rect 6040 65252 6096 65308
rect 6096 65252 6100 65308
rect 6036 65248 6100 65252
rect 36516 65308 36580 65312
rect 36516 65252 36520 65308
rect 36520 65252 36576 65308
rect 36576 65252 36580 65308
rect 36516 65248 36580 65252
rect 36596 65308 36660 65312
rect 36596 65252 36600 65308
rect 36600 65252 36656 65308
rect 36656 65252 36660 65308
rect 36596 65248 36660 65252
rect 36676 65308 36740 65312
rect 36676 65252 36680 65308
rect 36680 65252 36736 65308
rect 36736 65252 36740 65308
rect 36676 65248 36740 65252
rect 36756 65308 36820 65312
rect 36756 65252 36760 65308
rect 36760 65252 36816 65308
rect 36816 65252 36820 65308
rect 36756 65248 36820 65252
rect 67236 65308 67300 65312
rect 67236 65252 67240 65308
rect 67240 65252 67296 65308
rect 67296 65252 67300 65308
rect 67236 65248 67300 65252
rect 67316 65308 67380 65312
rect 67316 65252 67320 65308
rect 67320 65252 67376 65308
rect 67376 65252 67380 65308
rect 67316 65248 67380 65252
rect 67396 65308 67460 65312
rect 67396 65252 67400 65308
rect 67400 65252 67456 65308
rect 67456 65252 67460 65308
rect 67396 65248 67460 65252
rect 67476 65308 67540 65312
rect 67476 65252 67480 65308
rect 67480 65252 67536 65308
rect 67536 65252 67540 65308
rect 67476 65248 67540 65252
rect 5136 64764 5200 64768
rect 5136 64708 5140 64764
rect 5140 64708 5196 64764
rect 5196 64708 5200 64764
rect 5136 64704 5200 64708
rect 5216 64764 5280 64768
rect 5216 64708 5220 64764
rect 5220 64708 5276 64764
rect 5276 64708 5280 64764
rect 5216 64704 5280 64708
rect 5296 64764 5360 64768
rect 5296 64708 5300 64764
rect 5300 64708 5356 64764
rect 5356 64708 5360 64764
rect 5296 64704 5360 64708
rect 5376 64764 5440 64768
rect 5376 64708 5380 64764
rect 5380 64708 5436 64764
rect 5436 64708 5440 64764
rect 5376 64704 5440 64708
rect 35856 64764 35920 64768
rect 35856 64708 35860 64764
rect 35860 64708 35916 64764
rect 35916 64708 35920 64764
rect 35856 64704 35920 64708
rect 35936 64764 36000 64768
rect 35936 64708 35940 64764
rect 35940 64708 35996 64764
rect 35996 64708 36000 64764
rect 35936 64704 36000 64708
rect 36016 64764 36080 64768
rect 36016 64708 36020 64764
rect 36020 64708 36076 64764
rect 36076 64708 36080 64764
rect 36016 64704 36080 64708
rect 36096 64764 36160 64768
rect 36096 64708 36100 64764
rect 36100 64708 36156 64764
rect 36156 64708 36160 64764
rect 36096 64704 36160 64708
rect 66576 64764 66640 64768
rect 66576 64708 66580 64764
rect 66580 64708 66636 64764
rect 66636 64708 66640 64764
rect 66576 64704 66640 64708
rect 66656 64764 66720 64768
rect 66656 64708 66660 64764
rect 66660 64708 66716 64764
rect 66716 64708 66720 64764
rect 66656 64704 66720 64708
rect 66736 64764 66800 64768
rect 66736 64708 66740 64764
rect 66740 64708 66796 64764
rect 66796 64708 66800 64764
rect 66736 64704 66800 64708
rect 66816 64764 66880 64768
rect 66816 64708 66820 64764
rect 66820 64708 66876 64764
rect 66876 64708 66880 64764
rect 66816 64704 66880 64708
rect 5796 64220 5860 64224
rect 5796 64164 5800 64220
rect 5800 64164 5856 64220
rect 5856 64164 5860 64220
rect 5796 64160 5860 64164
rect 5876 64220 5940 64224
rect 5876 64164 5880 64220
rect 5880 64164 5936 64220
rect 5936 64164 5940 64220
rect 5876 64160 5940 64164
rect 5956 64220 6020 64224
rect 5956 64164 5960 64220
rect 5960 64164 6016 64220
rect 6016 64164 6020 64220
rect 5956 64160 6020 64164
rect 6036 64220 6100 64224
rect 6036 64164 6040 64220
rect 6040 64164 6096 64220
rect 6096 64164 6100 64220
rect 6036 64160 6100 64164
rect 36516 64220 36580 64224
rect 36516 64164 36520 64220
rect 36520 64164 36576 64220
rect 36576 64164 36580 64220
rect 36516 64160 36580 64164
rect 36596 64220 36660 64224
rect 36596 64164 36600 64220
rect 36600 64164 36656 64220
rect 36656 64164 36660 64220
rect 36596 64160 36660 64164
rect 36676 64220 36740 64224
rect 36676 64164 36680 64220
rect 36680 64164 36736 64220
rect 36736 64164 36740 64220
rect 36676 64160 36740 64164
rect 36756 64220 36820 64224
rect 36756 64164 36760 64220
rect 36760 64164 36816 64220
rect 36816 64164 36820 64220
rect 36756 64160 36820 64164
rect 67236 64220 67300 64224
rect 67236 64164 67240 64220
rect 67240 64164 67296 64220
rect 67296 64164 67300 64220
rect 67236 64160 67300 64164
rect 67316 64220 67380 64224
rect 67316 64164 67320 64220
rect 67320 64164 67376 64220
rect 67376 64164 67380 64220
rect 67316 64160 67380 64164
rect 67396 64220 67460 64224
rect 67396 64164 67400 64220
rect 67400 64164 67456 64220
rect 67456 64164 67460 64220
rect 67396 64160 67460 64164
rect 67476 64220 67540 64224
rect 67476 64164 67480 64220
rect 67480 64164 67536 64220
rect 67536 64164 67540 64220
rect 67476 64160 67540 64164
rect 5136 63676 5200 63680
rect 5136 63620 5140 63676
rect 5140 63620 5196 63676
rect 5196 63620 5200 63676
rect 5136 63616 5200 63620
rect 5216 63676 5280 63680
rect 5216 63620 5220 63676
rect 5220 63620 5276 63676
rect 5276 63620 5280 63676
rect 5216 63616 5280 63620
rect 5296 63676 5360 63680
rect 5296 63620 5300 63676
rect 5300 63620 5356 63676
rect 5356 63620 5360 63676
rect 5296 63616 5360 63620
rect 5376 63676 5440 63680
rect 5376 63620 5380 63676
rect 5380 63620 5436 63676
rect 5436 63620 5440 63676
rect 5376 63616 5440 63620
rect 35856 63676 35920 63680
rect 35856 63620 35860 63676
rect 35860 63620 35916 63676
rect 35916 63620 35920 63676
rect 35856 63616 35920 63620
rect 35936 63676 36000 63680
rect 35936 63620 35940 63676
rect 35940 63620 35996 63676
rect 35996 63620 36000 63676
rect 35936 63616 36000 63620
rect 36016 63676 36080 63680
rect 36016 63620 36020 63676
rect 36020 63620 36076 63676
rect 36076 63620 36080 63676
rect 36016 63616 36080 63620
rect 36096 63676 36160 63680
rect 36096 63620 36100 63676
rect 36100 63620 36156 63676
rect 36156 63620 36160 63676
rect 36096 63616 36160 63620
rect 66576 63676 66640 63680
rect 66576 63620 66580 63676
rect 66580 63620 66636 63676
rect 66636 63620 66640 63676
rect 66576 63616 66640 63620
rect 66656 63676 66720 63680
rect 66656 63620 66660 63676
rect 66660 63620 66716 63676
rect 66716 63620 66720 63676
rect 66656 63616 66720 63620
rect 66736 63676 66800 63680
rect 66736 63620 66740 63676
rect 66740 63620 66796 63676
rect 66796 63620 66800 63676
rect 66736 63616 66800 63620
rect 66816 63676 66880 63680
rect 66816 63620 66820 63676
rect 66820 63620 66876 63676
rect 66876 63620 66880 63676
rect 66816 63616 66880 63620
rect 5796 63132 5860 63136
rect 5796 63076 5800 63132
rect 5800 63076 5856 63132
rect 5856 63076 5860 63132
rect 5796 63072 5860 63076
rect 5876 63132 5940 63136
rect 5876 63076 5880 63132
rect 5880 63076 5936 63132
rect 5936 63076 5940 63132
rect 5876 63072 5940 63076
rect 5956 63132 6020 63136
rect 5956 63076 5960 63132
rect 5960 63076 6016 63132
rect 6016 63076 6020 63132
rect 5956 63072 6020 63076
rect 6036 63132 6100 63136
rect 6036 63076 6040 63132
rect 6040 63076 6096 63132
rect 6096 63076 6100 63132
rect 6036 63072 6100 63076
rect 36516 63132 36580 63136
rect 36516 63076 36520 63132
rect 36520 63076 36576 63132
rect 36576 63076 36580 63132
rect 36516 63072 36580 63076
rect 36596 63132 36660 63136
rect 36596 63076 36600 63132
rect 36600 63076 36656 63132
rect 36656 63076 36660 63132
rect 36596 63072 36660 63076
rect 36676 63132 36740 63136
rect 36676 63076 36680 63132
rect 36680 63076 36736 63132
rect 36736 63076 36740 63132
rect 36676 63072 36740 63076
rect 36756 63132 36820 63136
rect 36756 63076 36760 63132
rect 36760 63076 36816 63132
rect 36816 63076 36820 63132
rect 36756 63072 36820 63076
rect 67236 63132 67300 63136
rect 67236 63076 67240 63132
rect 67240 63076 67296 63132
rect 67296 63076 67300 63132
rect 67236 63072 67300 63076
rect 67316 63132 67380 63136
rect 67316 63076 67320 63132
rect 67320 63076 67376 63132
rect 67376 63076 67380 63132
rect 67316 63072 67380 63076
rect 67396 63132 67460 63136
rect 67396 63076 67400 63132
rect 67400 63076 67456 63132
rect 67456 63076 67460 63132
rect 67396 63072 67460 63076
rect 67476 63132 67540 63136
rect 67476 63076 67480 63132
rect 67480 63076 67536 63132
rect 67536 63076 67540 63132
rect 67476 63072 67540 63076
rect 5136 62588 5200 62592
rect 5136 62532 5140 62588
rect 5140 62532 5196 62588
rect 5196 62532 5200 62588
rect 5136 62528 5200 62532
rect 5216 62588 5280 62592
rect 5216 62532 5220 62588
rect 5220 62532 5276 62588
rect 5276 62532 5280 62588
rect 5216 62528 5280 62532
rect 5296 62588 5360 62592
rect 5296 62532 5300 62588
rect 5300 62532 5356 62588
rect 5356 62532 5360 62588
rect 5296 62528 5360 62532
rect 5376 62588 5440 62592
rect 5376 62532 5380 62588
rect 5380 62532 5436 62588
rect 5436 62532 5440 62588
rect 5376 62528 5440 62532
rect 35856 62588 35920 62592
rect 35856 62532 35860 62588
rect 35860 62532 35916 62588
rect 35916 62532 35920 62588
rect 35856 62528 35920 62532
rect 35936 62588 36000 62592
rect 35936 62532 35940 62588
rect 35940 62532 35996 62588
rect 35996 62532 36000 62588
rect 35936 62528 36000 62532
rect 36016 62588 36080 62592
rect 36016 62532 36020 62588
rect 36020 62532 36076 62588
rect 36076 62532 36080 62588
rect 36016 62528 36080 62532
rect 36096 62588 36160 62592
rect 36096 62532 36100 62588
rect 36100 62532 36156 62588
rect 36156 62532 36160 62588
rect 36096 62528 36160 62532
rect 66576 62588 66640 62592
rect 66576 62532 66580 62588
rect 66580 62532 66636 62588
rect 66636 62532 66640 62588
rect 66576 62528 66640 62532
rect 66656 62588 66720 62592
rect 66656 62532 66660 62588
rect 66660 62532 66716 62588
rect 66716 62532 66720 62588
rect 66656 62528 66720 62532
rect 66736 62588 66800 62592
rect 66736 62532 66740 62588
rect 66740 62532 66796 62588
rect 66796 62532 66800 62588
rect 66736 62528 66800 62532
rect 66816 62588 66880 62592
rect 66816 62532 66820 62588
rect 66820 62532 66876 62588
rect 66876 62532 66880 62588
rect 66816 62528 66880 62532
rect 5796 62044 5860 62048
rect 5796 61988 5800 62044
rect 5800 61988 5856 62044
rect 5856 61988 5860 62044
rect 5796 61984 5860 61988
rect 5876 62044 5940 62048
rect 5876 61988 5880 62044
rect 5880 61988 5936 62044
rect 5936 61988 5940 62044
rect 5876 61984 5940 61988
rect 5956 62044 6020 62048
rect 5956 61988 5960 62044
rect 5960 61988 6016 62044
rect 6016 61988 6020 62044
rect 5956 61984 6020 61988
rect 6036 62044 6100 62048
rect 6036 61988 6040 62044
rect 6040 61988 6096 62044
rect 6096 61988 6100 62044
rect 6036 61984 6100 61988
rect 36516 62044 36580 62048
rect 36516 61988 36520 62044
rect 36520 61988 36576 62044
rect 36576 61988 36580 62044
rect 36516 61984 36580 61988
rect 36596 62044 36660 62048
rect 36596 61988 36600 62044
rect 36600 61988 36656 62044
rect 36656 61988 36660 62044
rect 36596 61984 36660 61988
rect 36676 62044 36740 62048
rect 36676 61988 36680 62044
rect 36680 61988 36736 62044
rect 36736 61988 36740 62044
rect 36676 61984 36740 61988
rect 36756 62044 36820 62048
rect 36756 61988 36760 62044
rect 36760 61988 36816 62044
rect 36816 61988 36820 62044
rect 36756 61984 36820 61988
rect 67236 62044 67300 62048
rect 67236 61988 67240 62044
rect 67240 61988 67296 62044
rect 67296 61988 67300 62044
rect 67236 61984 67300 61988
rect 67316 62044 67380 62048
rect 67316 61988 67320 62044
rect 67320 61988 67376 62044
rect 67376 61988 67380 62044
rect 67316 61984 67380 61988
rect 67396 62044 67460 62048
rect 67396 61988 67400 62044
rect 67400 61988 67456 62044
rect 67456 61988 67460 62044
rect 67396 61984 67460 61988
rect 67476 62044 67540 62048
rect 67476 61988 67480 62044
rect 67480 61988 67536 62044
rect 67536 61988 67540 62044
rect 67476 61984 67540 61988
rect 5136 61500 5200 61504
rect 5136 61444 5140 61500
rect 5140 61444 5196 61500
rect 5196 61444 5200 61500
rect 5136 61440 5200 61444
rect 5216 61500 5280 61504
rect 5216 61444 5220 61500
rect 5220 61444 5276 61500
rect 5276 61444 5280 61500
rect 5216 61440 5280 61444
rect 5296 61500 5360 61504
rect 5296 61444 5300 61500
rect 5300 61444 5356 61500
rect 5356 61444 5360 61500
rect 5296 61440 5360 61444
rect 5376 61500 5440 61504
rect 5376 61444 5380 61500
rect 5380 61444 5436 61500
rect 5436 61444 5440 61500
rect 5376 61440 5440 61444
rect 35856 61500 35920 61504
rect 35856 61444 35860 61500
rect 35860 61444 35916 61500
rect 35916 61444 35920 61500
rect 35856 61440 35920 61444
rect 35936 61500 36000 61504
rect 35936 61444 35940 61500
rect 35940 61444 35996 61500
rect 35996 61444 36000 61500
rect 35936 61440 36000 61444
rect 36016 61500 36080 61504
rect 36016 61444 36020 61500
rect 36020 61444 36076 61500
rect 36076 61444 36080 61500
rect 36016 61440 36080 61444
rect 36096 61500 36160 61504
rect 36096 61444 36100 61500
rect 36100 61444 36156 61500
rect 36156 61444 36160 61500
rect 36096 61440 36160 61444
rect 66576 61500 66640 61504
rect 66576 61444 66580 61500
rect 66580 61444 66636 61500
rect 66636 61444 66640 61500
rect 66576 61440 66640 61444
rect 66656 61500 66720 61504
rect 66656 61444 66660 61500
rect 66660 61444 66716 61500
rect 66716 61444 66720 61500
rect 66656 61440 66720 61444
rect 66736 61500 66800 61504
rect 66736 61444 66740 61500
rect 66740 61444 66796 61500
rect 66796 61444 66800 61500
rect 66736 61440 66800 61444
rect 66816 61500 66880 61504
rect 66816 61444 66820 61500
rect 66820 61444 66876 61500
rect 66876 61444 66880 61500
rect 66816 61440 66880 61444
rect 5796 60956 5860 60960
rect 5796 60900 5800 60956
rect 5800 60900 5856 60956
rect 5856 60900 5860 60956
rect 5796 60896 5860 60900
rect 5876 60956 5940 60960
rect 5876 60900 5880 60956
rect 5880 60900 5936 60956
rect 5936 60900 5940 60956
rect 5876 60896 5940 60900
rect 5956 60956 6020 60960
rect 5956 60900 5960 60956
rect 5960 60900 6016 60956
rect 6016 60900 6020 60956
rect 5956 60896 6020 60900
rect 6036 60956 6100 60960
rect 6036 60900 6040 60956
rect 6040 60900 6096 60956
rect 6096 60900 6100 60956
rect 6036 60896 6100 60900
rect 36516 60956 36580 60960
rect 36516 60900 36520 60956
rect 36520 60900 36576 60956
rect 36576 60900 36580 60956
rect 36516 60896 36580 60900
rect 36596 60956 36660 60960
rect 36596 60900 36600 60956
rect 36600 60900 36656 60956
rect 36656 60900 36660 60956
rect 36596 60896 36660 60900
rect 36676 60956 36740 60960
rect 36676 60900 36680 60956
rect 36680 60900 36736 60956
rect 36736 60900 36740 60956
rect 36676 60896 36740 60900
rect 36756 60956 36820 60960
rect 36756 60900 36760 60956
rect 36760 60900 36816 60956
rect 36816 60900 36820 60956
rect 36756 60896 36820 60900
rect 67236 60956 67300 60960
rect 67236 60900 67240 60956
rect 67240 60900 67296 60956
rect 67296 60900 67300 60956
rect 67236 60896 67300 60900
rect 67316 60956 67380 60960
rect 67316 60900 67320 60956
rect 67320 60900 67376 60956
rect 67376 60900 67380 60956
rect 67316 60896 67380 60900
rect 67396 60956 67460 60960
rect 67396 60900 67400 60956
rect 67400 60900 67456 60956
rect 67456 60900 67460 60956
rect 67396 60896 67460 60900
rect 67476 60956 67540 60960
rect 67476 60900 67480 60956
rect 67480 60900 67536 60956
rect 67536 60900 67540 60956
rect 67476 60896 67540 60900
rect 5136 60412 5200 60416
rect 5136 60356 5140 60412
rect 5140 60356 5196 60412
rect 5196 60356 5200 60412
rect 5136 60352 5200 60356
rect 5216 60412 5280 60416
rect 5216 60356 5220 60412
rect 5220 60356 5276 60412
rect 5276 60356 5280 60412
rect 5216 60352 5280 60356
rect 5296 60412 5360 60416
rect 5296 60356 5300 60412
rect 5300 60356 5356 60412
rect 5356 60356 5360 60412
rect 5296 60352 5360 60356
rect 5376 60412 5440 60416
rect 5376 60356 5380 60412
rect 5380 60356 5436 60412
rect 5436 60356 5440 60412
rect 5376 60352 5440 60356
rect 35856 60412 35920 60416
rect 35856 60356 35860 60412
rect 35860 60356 35916 60412
rect 35916 60356 35920 60412
rect 35856 60352 35920 60356
rect 35936 60412 36000 60416
rect 35936 60356 35940 60412
rect 35940 60356 35996 60412
rect 35996 60356 36000 60412
rect 35936 60352 36000 60356
rect 36016 60412 36080 60416
rect 36016 60356 36020 60412
rect 36020 60356 36076 60412
rect 36076 60356 36080 60412
rect 36016 60352 36080 60356
rect 36096 60412 36160 60416
rect 36096 60356 36100 60412
rect 36100 60356 36156 60412
rect 36156 60356 36160 60412
rect 36096 60352 36160 60356
rect 66576 60412 66640 60416
rect 66576 60356 66580 60412
rect 66580 60356 66636 60412
rect 66636 60356 66640 60412
rect 66576 60352 66640 60356
rect 66656 60412 66720 60416
rect 66656 60356 66660 60412
rect 66660 60356 66716 60412
rect 66716 60356 66720 60412
rect 66656 60352 66720 60356
rect 66736 60412 66800 60416
rect 66736 60356 66740 60412
rect 66740 60356 66796 60412
rect 66796 60356 66800 60412
rect 66736 60352 66800 60356
rect 66816 60412 66880 60416
rect 66816 60356 66820 60412
rect 66820 60356 66876 60412
rect 66876 60356 66880 60412
rect 66816 60352 66880 60356
rect 5796 59868 5860 59872
rect 5796 59812 5800 59868
rect 5800 59812 5856 59868
rect 5856 59812 5860 59868
rect 5796 59808 5860 59812
rect 5876 59868 5940 59872
rect 5876 59812 5880 59868
rect 5880 59812 5936 59868
rect 5936 59812 5940 59868
rect 5876 59808 5940 59812
rect 5956 59868 6020 59872
rect 5956 59812 5960 59868
rect 5960 59812 6016 59868
rect 6016 59812 6020 59868
rect 5956 59808 6020 59812
rect 6036 59868 6100 59872
rect 6036 59812 6040 59868
rect 6040 59812 6096 59868
rect 6096 59812 6100 59868
rect 6036 59808 6100 59812
rect 36516 59868 36580 59872
rect 36516 59812 36520 59868
rect 36520 59812 36576 59868
rect 36576 59812 36580 59868
rect 36516 59808 36580 59812
rect 36596 59868 36660 59872
rect 36596 59812 36600 59868
rect 36600 59812 36656 59868
rect 36656 59812 36660 59868
rect 36596 59808 36660 59812
rect 36676 59868 36740 59872
rect 36676 59812 36680 59868
rect 36680 59812 36736 59868
rect 36736 59812 36740 59868
rect 36676 59808 36740 59812
rect 36756 59868 36820 59872
rect 36756 59812 36760 59868
rect 36760 59812 36816 59868
rect 36816 59812 36820 59868
rect 36756 59808 36820 59812
rect 67236 59868 67300 59872
rect 67236 59812 67240 59868
rect 67240 59812 67296 59868
rect 67296 59812 67300 59868
rect 67236 59808 67300 59812
rect 67316 59868 67380 59872
rect 67316 59812 67320 59868
rect 67320 59812 67376 59868
rect 67376 59812 67380 59868
rect 67316 59808 67380 59812
rect 67396 59868 67460 59872
rect 67396 59812 67400 59868
rect 67400 59812 67456 59868
rect 67456 59812 67460 59868
rect 67396 59808 67460 59812
rect 67476 59868 67540 59872
rect 67476 59812 67480 59868
rect 67480 59812 67536 59868
rect 67536 59812 67540 59868
rect 67476 59808 67540 59812
rect 5136 59324 5200 59328
rect 5136 59268 5140 59324
rect 5140 59268 5196 59324
rect 5196 59268 5200 59324
rect 5136 59264 5200 59268
rect 5216 59324 5280 59328
rect 5216 59268 5220 59324
rect 5220 59268 5276 59324
rect 5276 59268 5280 59324
rect 5216 59264 5280 59268
rect 5296 59324 5360 59328
rect 5296 59268 5300 59324
rect 5300 59268 5356 59324
rect 5356 59268 5360 59324
rect 5296 59264 5360 59268
rect 5376 59324 5440 59328
rect 5376 59268 5380 59324
rect 5380 59268 5436 59324
rect 5436 59268 5440 59324
rect 5376 59264 5440 59268
rect 35856 59324 35920 59328
rect 35856 59268 35860 59324
rect 35860 59268 35916 59324
rect 35916 59268 35920 59324
rect 35856 59264 35920 59268
rect 35936 59324 36000 59328
rect 35936 59268 35940 59324
rect 35940 59268 35996 59324
rect 35996 59268 36000 59324
rect 35936 59264 36000 59268
rect 36016 59324 36080 59328
rect 36016 59268 36020 59324
rect 36020 59268 36076 59324
rect 36076 59268 36080 59324
rect 36016 59264 36080 59268
rect 36096 59324 36160 59328
rect 36096 59268 36100 59324
rect 36100 59268 36156 59324
rect 36156 59268 36160 59324
rect 36096 59264 36160 59268
rect 66576 59324 66640 59328
rect 66576 59268 66580 59324
rect 66580 59268 66636 59324
rect 66636 59268 66640 59324
rect 66576 59264 66640 59268
rect 66656 59324 66720 59328
rect 66656 59268 66660 59324
rect 66660 59268 66716 59324
rect 66716 59268 66720 59324
rect 66656 59264 66720 59268
rect 66736 59324 66800 59328
rect 66736 59268 66740 59324
rect 66740 59268 66796 59324
rect 66796 59268 66800 59324
rect 66736 59264 66800 59268
rect 66816 59324 66880 59328
rect 66816 59268 66820 59324
rect 66820 59268 66876 59324
rect 66876 59268 66880 59324
rect 66816 59264 66880 59268
rect 5796 58780 5860 58784
rect 5796 58724 5800 58780
rect 5800 58724 5856 58780
rect 5856 58724 5860 58780
rect 5796 58720 5860 58724
rect 5876 58780 5940 58784
rect 5876 58724 5880 58780
rect 5880 58724 5936 58780
rect 5936 58724 5940 58780
rect 5876 58720 5940 58724
rect 5956 58780 6020 58784
rect 5956 58724 5960 58780
rect 5960 58724 6016 58780
rect 6016 58724 6020 58780
rect 5956 58720 6020 58724
rect 6036 58780 6100 58784
rect 6036 58724 6040 58780
rect 6040 58724 6096 58780
rect 6096 58724 6100 58780
rect 6036 58720 6100 58724
rect 36516 58780 36580 58784
rect 36516 58724 36520 58780
rect 36520 58724 36576 58780
rect 36576 58724 36580 58780
rect 36516 58720 36580 58724
rect 36596 58780 36660 58784
rect 36596 58724 36600 58780
rect 36600 58724 36656 58780
rect 36656 58724 36660 58780
rect 36596 58720 36660 58724
rect 36676 58780 36740 58784
rect 36676 58724 36680 58780
rect 36680 58724 36736 58780
rect 36736 58724 36740 58780
rect 36676 58720 36740 58724
rect 36756 58780 36820 58784
rect 36756 58724 36760 58780
rect 36760 58724 36816 58780
rect 36816 58724 36820 58780
rect 36756 58720 36820 58724
rect 67236 58780 67300 58784
rect 67236 58724 67240 58780
rect 67240 58724 67296 58780
rect 67296 58724 67300 58780
rect 67236 58720 67300 58724
rect 67316 58780 67380 58784
rect 67316 58724 67320 58780
rect 67320 58724 67376 58780
rect 67376 58724 67380 58780
rect 67316 58720 67380 58724
rect 67396 58780 67460 58784
rect 67396 58724 67400 58780
rect 67400 58724 67456 58780
rect 67456 58724 67460 58780
rect 67396 58720 67460 58724
rect 67476 58780 67540 58784
rect 67476 58724 67480 58780
rect 67480 58724 67536 58780
rect 67536 58724 67540 58780
rect 67476 58720 67540 58724
rect 5136 58236 5200 58240
rect 5136 58180 5140 58236
rect 5140 58180 5196 58236
rect 5196 58180 5200 58236
rect 5136 58176 5200 58180
rect 5216 58236 5280 58240
rect 5216 58180 5220 58236
rect 5220 58180 5276 58236
rect 5276 58180 5280 58236
rect 5216 58176 5280 58180
rect 5296 58236 5360 58240
rect 5296 58180 5300 58236
rect 5300 58180 5356 58236
rect 5356 58180 5360 58236
rect 5296 58176 5360 58180
rect 5376 58236 5440 58240
rect 5376 58180 5380 58236
rect 5380 58180 5436 58236
rect 5436 58180 5440 58236
rect 5376 58176 5440 58180
rect 35856 58236 35920 58240
rect 35856 58180 35860 58236
rect 35860 58180 35916 58236
rect 35916 58180 35920 58236
rect 35856 58176 35920 58180
rect 35936 58236 36000 58240
rect 35936 58180 35940 58236
rect 35940 58180 35996 58236
rect 35996 58180 36000 58236
rect 35936 58176 36000 58180
rect 36016 58236 36080 58240
rect 36016 58180 36020 58236
rect 36020 58180 36076 58236
rect 36076 58180 36080 58236
rect 36016 58176 36080 58180
rect 36096 58236 36160 58240
rect 36096 58180 36100 58236
rect 36100 58180 36156 58236
rect 36156 58180 36160 58236
rect 36096 58176 36160 58180
rect 66576 58236 66640 58240
rect 66576 58180 66580 58236
rect 66580 58180 66636 58236
rect 66636 58180 66640 58236
rect 66576 58176 66640 58180
rect 66656 58236 66720 58240
rect 66656 58180 66660 58236
rect 66660 58180 66716 58236
rect 66716 58180 66720 58236
rect 66656 58176 66720 58180
rect 66736 58236 66800 58240
rect 66736 58180 66740 58236
rect 66740 58180 66796 58236
rect 66796 58180 66800 58236
rect 66736 58176 66800 58180
rect 66816 58236 66880 58240
rect 66816 58180 66820 58236
rect 66820 58180 66876 58236
rect 66876 58180 66880 58236
rect 66816 58176 66880 58180
rect 5796 57692 5860 57696
rect 5796 57636 5800 57692
rect 5800 57636 5856 57692
rect 5856 57636 5860 57692
rect 5796 57632 5860 57636
rect 5876 57692 5940 57696
rect 5876 57636 5880 57692
rect 5880 57636 5936 57692
rect 5936 57636 5940 57692
rect 5876 57632 5940 57636
rect 5956 57692 6020 57696
rect 5956 57636 5960 57692
rect 5960 57636 6016 57692
rect 6016 57636 6020 57692
rect 5956 57632 6020 57636
rect 6036 57692 6100 57696
rect 6036 57636 6040 57692
rect 6040 57636 6096 57692
rect 6096 57636 6100 57692
rect 6036 57632 6100 57636
rect 36516 57692 36580 57696
rect 36516 57636 36520 57692
rect 36520 57636 36576 57692
rect 36576 57636 36580 57692
rect 36516 57632 36580 57636
rect 36596 57692 36660 57696
rect 36596 57636 36600 57692
rect 36600 57636 36656 57692
rect 36656 57636 36660 57692
rect 36596 57632 36660 57636
rect 36676 57692 36740 57696
rect 36676 57636 36680 57692
rect 36680 57636 36736 57692
rect 36736 57636 36740 57692
rect 36676 57632 36740 57636
rect 36756 57692 36820 57696
rect 36756 57636 36760 57692
rect 36760 57636 36816 57692
rect 36816 57636 36820 57692
rect 36756 57632 36820 57636
rect 67236 57692 67300 57696
rect 67236 57636 67240 57692
rect 67240 57636 67296 57692
rect 67296 57636 67300 57692
rect 67236 57632 67300 57636
rect 67316 57692 67380 57696
rect 67316 57636 67320 57692
rect 67320 57636 67376 57692
rect 67376 57636 67380 57692
rect 67316 57632 67380 57636
rect 67396 57692 67460 57696
rect 67396 57636 67400 57692
rect 67400 57636 67456 57692
rect 67456 57636 67460 57692
rect 67396 57632 67460 57636
rect 67476 57692 67540 57696
rect 67476 57636 67480 57692
rect 67480 57636 67536 57692
rect 67536 57636 67540 57692
rect 67476 57632 67540 57636
rect 5136 57148 5200 57152
rect 5136 57092 5140 57148
rect 5140 57092 5196 57148
rect 5196 57092 5200 57148
rect 5136 57088 5200 57092
rect 5216 57148 5280 57152
rect 5216 57092 5220 57148
rect 5220 57092 5276 57148
rect 5276 57092 5280 57148
rect 5216 57088 5280 57092
rect 5296 57148 5360 57152
rect 5296 57092 5300 57148
rect 5300 57092 5356 57148
rect 5356 57092 5360 57148
rect 5296 57088 5360 57092
rect 5376 57148 5440 57152
rect 5376 57092 5380 57148
rect 5380 57092 5436 57148
rect 5436 57092 5440 57148
rect 5376 57088 5440 57092
rect 35856 57148 35920 57152
rect 35856 57092 35860 57148
rect 35860 57092 35916 57148
rect 35916 57092 35920 57148
rect 35856 57088 35920 57092
rect 35936 57148 36000 57152
rect 35936 57092 35940 57148
rect 35940 57092 35996 57148
rect 35996 57092 36000 57148
rect 35936 57088 36000 57092
rect 36016 57148 36080 57152
rect 36016 57092 36020 57148
rect 36020 57092 36076 57148
rect 36076 57092 36080 57148
rect 36016 57088 36080 57092
rect 36096 57148 36160 57152
rect 36096 57092 36100 57148
rect 36100 57092 36156 57148
rect 36156 57092 36160 57148
rect 36096 57088 36160 57092
rect 66576 57148 66640 57152
rect 66576 57092 66580 57148
rect 66580 57092 66636 57148
rect 66636 57092 66640 57148
rect 66576 57088 66640 57092
rect 66656 57148 66720 57152
rect 66656 57092 66660 57148
rect 66660 57092 66716 57148
rect 66716 57092 66720 57148
rect 66656 57088 66720 57092
rect 66736 57148 66800 57152
rect 66736 57092 66740 57148
rect 66740 57092 66796 57148
rect 66796 57092 66800 57148
rect 66736 57088 66800 57092
rect 66816 57148 66880 57152
rect 66816 57092 66820 57148
rect 66820 57092 66876 57148
rect 66876 57092 66880 57148
rect 66816 57088 66880 57092
rect 5796 56604 5860 56608
rect 5796 56548 5800 56604
rect 5800 56548 5856 56604
rect 5856 56548 5860 56604
rect 5796 56544 5860 56548
rect 5876 56604 5940 56608
rect 5876 56548 5880 56604
rect 5880 56548 5936 56604
rect 5936 56548 5940 56604
rect 5876 56544 5940 56548
rect 5956 56604 6020 56608
rect 5956 56548 5960 56604
rect 5960 56548 6016 56604
rect 6016 56548 6020 56604
rect 5956 56544 6020 56548
rect 6036 56604 6100 56608
rect 6036 56548 6040 56604
rect 6040 56548 6096 56604
rect 6096 56548 6100 56604
rect 6036 56544 6100 56548
rect 36516 56604 36580 56608
rect 36516 56548 36520 56604
rect 36520 56548 36576 56604
rect 36576 56548 36580 56604
rect 36516 56544 36580 56548
rect 36596 56604 36660 56608
rect 36596 56548 36600 56604
rect 36600 56548 36656 56604
rect 36656 56548 36660 56604
rect 36596 56544 36660 56548
rect 36676 56604 36740 56608
rect 36676 56548 36680 56604
rect 36680 56548 36736 56604
rect 36736 56548 36740 56604
rect 36676 56544 36740 56548
rect 36756 56604 36820 56608
rect 36756 56548 36760 56604
rect 36760 56548 36816 56604
rect 36816 56548 36820 56604
rect 36756 56544 36820 56548
rect 67236 56604 67300 56608
rect 67236 56548 67240 56604
rect 67240 56548 67296 56604
rect 67296 56548 67300 56604
rect 67236 56544 67300 56548
rect 67316 56604 67380 56608
rect 67316 56548 67320 56604
rect 67320 56548 67376 56604
rect 67376 56548 67380 56604
rect 67316 56544 67380 56548
rect 67396 56604 67460 56608
rect 67396 56548 67400 56604
rect 67400 56548 67456 56604
rect 67456 56548 67460 56604
rect 67396 56544 67460 56548
rect 67476 56604 67540 56608
rect 67476 56548 67480 56604
rect 67480 56548 67536 56604
rect 67536 56548 67540 56604
rect 67476 56544 67540 56548
rect 5136 56060 5200 56064
rect 5136 56004 5140 56060
rect 5140 56004 5196 56060
rect 5196 56004 5200 56060
rect 5136 56000 5200 56004
rect 5216 56060 5280 56064
rect 5216 56004 5220 56060
rect 5220 56004 5276 56060
rect 5276 56004 5280 56060
rect 5216 56000 5280 56004
rect 5296 56060 5360 56064
rect 5296 56004 5300 56060
rect 5300 56004 5356 56060
rect 5356 56004 5360 56060
rect 5296 56000 5360 56004
rect 5376 56060 5440 56064
rect 5376 56004 5380 56060
rect 5380 56004 5436 56060
rect 5436 56004 5440 56060
rect 5376 56000 5440 56004
rect 35856 56060 35920 56064
rect 35856 56004 35860 56060
rect 35860 56004 35916 56060
rect 35916 56004 35920 56060
rect 35856 56000 35920 56004
rect 35936 56060 36000 56064
rect 35936 56004 35940 56060
rect 35940 56004 35996 56060
rect 35996 56004 36000 56060
rect 35936 56000 36000 56004
rect 36016 56060 36080 56064
rect 36016 56004 36020 56060
rect 36020 56004 36076 56060
rect 36076 56004 36080 56060
rect 36016 56000 36080 56004
rect 36096 56060 36160 56064
rect 36096 56004 36100 56060
rect 36100 56004 36156 56060
rect 36156 56004 36160 56060
rect 36096 56000 36160 56004
rect 66576 56060 66640 56064
rect 66576 56004 66580 56060
rect 66580 56004 66636 56060
rect 66636 56004 66640 56060
rect 66576 56000 66640 56004
rect 66656 56060 66720 56064
rect 66656 56004 66660 56060
rect 66660 56004 66716 56060
rect 66716 56004 66720 56060
rect 66656 56000 66720 56004
rect 66736 56060 66800 56064
rect 66736 56004 66740 56060
rect 66740 56004 66796 56060
rect 66796 56004 66800 56060
rect 66736 56000 66800 56004
rect 66816 56060 66880 56064
rect 66816 56004 66820 56060
rect 66820 56004 66876 56060
rect 66876 56004 66880 56060
rect 66816 56000 66880 56004
rect 5796 55516 5860 55520
rect 5796 55460 5800 55516
rect 5800 55460 5856 55516
rect 5856 55460 5860 55516
rect 5796 55456 5860 55460
rect 5876 55516 5940 55520
rect 5876 55460 5880 55516
rect 5880 55460 5936 55516
rect 5936 55460 5940 55516
rect 5876 55456 5940 55460
rect 5956 55516 6020 55520
rect 5956 55460 5960 55516
rect 5960 55460 6016 55516
rect 6016 55460 6020 55516
rect 5956 55456 6020 55460
rect 6036 55516 6100 55520
rect 6036 55460 6040 55516
rect 6040 55460 6096 55516
rect 6096 55460 6100 55516
rect 6036 55456 6100 55460
rect 36516 55516 36580 55520
rect 36516 55460 36520 55516
rect 36520 55460 36576 55516
rect 36576 55460 36580 55516
rect 36516 55456 36580 55460
rect 36596 55516 36660 55520
rect 36596 55460 36600 55516
rect 36600 55460 36656 55516
rect 36656 55460 36660 55516
rect 36596 55456 36660 55460
rect 36676 55516 36740 55520
rect 36676 55460 36680 55516
rect 36680 55460 36736 55516
rect 36736 55460 36740 55516
rect 36676 55456 36740 55460
rect 36756 55516 36820 55520
rect 36756 55460 36760 55516
rect 36760 55460 36816 55516
rect 36816 55460 36820 55516
rect 36756 55456 36820 55460
rect 67236 55516 67300 55520
rect 67236 55460 67240 55516
rect 67240 55460 67296 55516
rect 67296 55460 67300 55516
rect 67236 55456 67300 55460
rect 67316 55516 67380 55520
rect 67316 55460 67320 55516
rect 67320 55460 67376 55516
rect 67376 55460 67380 55516
rect 67316 55456 67380 55460
rect 67396 55516 67460 55520
rect 67396 55460 67400 55516
rect 67400 55460 67456 55516
rect 67456 55460 67460 55516
rect 67396 55456 67460 55460
rect 67476 55516 67540 55520
rect 67476 55460 67480 55516
rect 67480 55460 67536 55516
rect 67536 55460 67540 55516
rect 67476 55456 67540 55460
rect 5136 54972 5200 54976
rect 5136 54916 5140 54972
rect 5140 54916 5196 54972
rect 5196 54916 5200 54972
rect 5136 54912 5200 54916
rect 5216 54972 5280 54976
rect 5216 54916 5220 54972
rect 5220 54916 5276 54972
rect 5276 54916 5280 54972
rect 5216 54912 5280 54916
rect 5296 54972 5360 54976
rect 5296 54916 5300 54972
rect 5300 54916 5356 54972
rect 5356 54916 5360 54972
rect 5296 54912 5360 54916
rect 5376 54972 5440 54976
rect 5376 54916 5380 54972
rect 5380 54916 5436 54972
rect 5436 54916 5440 54972
rect 5376 54912 5440 54916
rect 35856 54972 35920 54976
rect 35856 54916 35860 54972
rect 35860 54916 35916 54972
rect 35916 54916 35920 54972
rect 35856 54912 35920 54916
rect 35936 54972 36000 54976
rect 35936 54916 35940 54972
rect 35940 54916 35996 54972
rect 35996 54916 36000 54972
rect 35936 54912 36000 54916
rect 36016 54972 36080 54976
rect 36016 54916 36020 54972
rect 36020 54916 36076 54972
rect 36076 54916 36080 54972
rect 36016 54912 36080 54916
rect 36096 54972 36160 54976
rect 36096 54916 36100 54972
rect 36100 54916 36156 54972
rect 36156 54916 36160 54972
rect 36096 54912 36160 54916
rect 66576 54972 66640 54976
rect 66576 54916 66580 54972
rect 66580 54916 66636 54972
rect 66636 54916 66640 54972
rect 66576 54912 66640 54916
rect 66656 54972 66720 54976
rect 66656 54916 66660 54972
rect 66660 54916 66716 54972
rect 66716 54916 66720 54972
rect 66656 54912 66720 54916
rect 66736 54972 66800 54976
rect 66736 54916 66740 54972
rect 66740 54916 66796 54972
rect 66796 54916 66800 54972
rect 66736 54912 66800 54916
rect 66816 54972 66880 54976
rect 66816 54916 66820 54972
rect 66820 54916 66876 54972
rect 66876 54916 66880 54972
rect 66816 54912 66880 54916
rect 5796 54428 5860 54432
rect 5796 54372 5800 54428
rect 5800 54372 5856 54428
rect 5856 54372 5860 54428
rect 5796 54368 5860 54372
rect 5876 54428 5940 54432
rect 5876 54372 5880 54428
rect 5880 54372 5936 54428
rect 5936 54372 5940 54428
rect 5876 54368 5940 54372
rect 5956 54428 6020 54432
rect 5956 54372 5960 54428
rect 5960 54372 6016 54428
rect 6016 54372 6020 54428
rect 5956 54368 6020 54372
rect 6036 54428 6100 54432
rect 6036 54372 6040 54428
rect 6040 54372 6096 54428
rect 6096 54372 6100 54428
rect 6036 54368 6100 54372
rect 36516 54428 36580 54432
rect 36516 54372 36520 54428
rect 36520 54372 36576 54428
rect 36576 54372 36580 54428
rect 36516 54368 36580 54372
rect 36596 54428 36660 54432
rect 36596 54372 36600 54428
rect 36600 54372 36656 54428
rect 36656 54372 36660 54428
rect 36596 54368 36660 54372
rect 36676 54428 36740 54432
rect 36676 54372 36680 54428
rect 36680 54372 36736 54428
rect 36736 54372 36740 54428
rect 36676 54368 36740 54372
rect 36756 54428 36820 54432
rect 36756 54372 36760 54428
rect 36760 54372 36816 54428
rect 36816 54372 36820 54428
rect 36756 54368 36820 54372
rect 67236 54428 67300 54432
rect 67236 54372 67240 54428
rect 67240 54372 67296 54428
rect 67296 54372 67300 54428
rect 67236 54368 67300 54372
rect 67316 54428 67380 54432
rect 67316 54372 67320 54428
rect 67320 54372 67376 54428
rect 67376 54372 67380 54428
rect 67316 54368 67380 54372
rect 67396 54428 67460 54432
rect 67396 54372 67400 54428
rect 67400 54372 67456 54428
rect 67456 54372 67460 54428
rect 67396 54368 67460 54372
rect 67476 54428 67540 54432
rect 67476 54372 67480 54428
rect 67480 54372 67536 54428
rect 67536 54372 67540 54428
rect 67476 54368 67540 54372
rect 5136 53884 5200 53888
rect 5136 53828 5140 53884
rect 5140 53828 5196 53884
rect 5196 53828 5200 53884
rect 5136 53824 5200 53828
rect 5216 53884 5280 53888
rect 5216 53828 5220 53884
rect 5220 53828 5276 53884
rect 5276 53828 5280 53884
rect 5216 53824 5280 53828
rect 5296 53884 5360 53888
rect 5296 53828 5300 53884
rect 5300 53828 5356 53884
rect 5356 53828 5360 53884
rect 5296 53824 5360 53828
rect 5376 53884 5440 53888
rect 5376 53828 5380 53884
rect 5380 53828 5436 53884
rect 5436 53828 5440 53884
rect 5376 53824 5440 53828
rect 35856 53884 35920 53888
rect 35856 53828 35860 53884
rect 35860 53828 35916 53884
rect 35916 53828 35920 53884
rect 35856 53824 35920 53828
rect 35936 53884 36000 53888
rect 35936 53828 35940 53884
rect 35940 53828 35996 53884
rect 35996 53828 36000 53884
rect 35936 53824 36000 53828
rect 36016 53884 36080 53888
rect 36016 53828 36020 53884
rect 36020 53828 36076 53884
rect 36076 53828 36080 53884
rect 36016 53824 36080 53828
rect 36096 53884 36160 53888
rect 36096 53828 36100 53884
rect 36100 53828 36156 53884
rect 36156 53828 36160 53884
rect 36096 53824 36160 53828
rect 66576 53884 66640 53888
rect 66576 53828 66580 53884
rect 66580 53828 66636 53884
rect 66636 53828 66640 53884
rect 66576 53824 66640 53828
rect 66656 53884 66720 53888
rect 66656 53828 66660 53884
rect 66660 53828 66716 53884
rect 66716 53828 66720 53884
rect 66656 53824 66720 53828
rect 66736 53884 66800 53888
rect 66736 53828 66740 53884
rect 66740 53828 66796 53884
rect 66796 53828 66800 53884
rect 66736 53824 66800 53828
rect 66816 53884 66880 53888
rect 66816 53828 66820 53884
rect 66820 53828 66876 53884
rect 66876 53828 66880 53884
rect 66816 53824 66880 53828
rect 5796 53340 5860 53344
rect 5796 53284 5800 53340
rect 5800 53284 5856 53340
rect 5856 53284 5860 53340
rect 5796 53280 5860 53284
rect 5876 53340 5940 53344
rect 5876 53284 5880 53340
rect 5880 53284 5936 53340
rect 5936 53284 5940 53340
rect 5876 53280 5940 53284
rect 5956 53340 6020 53344
rect 5956 53284 5960 53340
rect 5960 53284 6016 53340
rect 6016 53284 6020 53340
rect 5956 53280 6020 53284
rect 6036 53340 6100 53344
rect 6036 53284 6040 53340
rect 6040 53284 6096 53340
rect 6096 53284 6100 53340
rect 6036 53280 6100 53284
rect 36516 53340 36580 53344
rect 36516 53284 36520 53340
rect 36520 53284 36576 53340
rect 36576 53284 36580 53340
rect 36516 53280 36580 53284
rect 36596 53340 36660 53344
rect 36596 53284 36600 53340
rect 36600 53284 36656 53340
rect 36656 53284 36660 53340
rect 36596 53280 36660 53284
rect 36676 53340 36740 53344
rect 36676 53284 36680 53340
rect 36680 53284 36736 53340
rect 36736 53284 36740 53340
rect 36676 53280 36740 53284
rect 36756 53340 36820 53344
rect 36756 53284 36760 53340
rect 36760 53284 36816 53340
rect 36816 53284 36820 53340
rect 36756 53280 36820 53284
rect 67236 53340 67300 53344
rect 67236 53284 67240 53340
rect 67240 53284 67296 53340
rect 67296 53284 67300 53340
rect 67236 53280 67300 53284
rect 67316 53340 67380 53344
rect 67316 53284 67320 53340
rect 67320 53284 67376 53340
rect 67376 53284 67380 53340
rect 67316 53280 67380 53284
rect 67396 53340 67460 53344
rect 67396 53284 67400 53340
rect 67400 53284 67456 53340
rect 67456 53284 67460 53340
rect 67396 53280 67460 53284
rect 67476 53340 67540 53344
rect 67476 53284 67480 53340
rect 67480 53284 67536 53340
rect 67536 53284 67540 53340
rect 67476 53280 67540 53284
rect 5136 52796 5200 52800
rect 5136 52740 5140 52796
rect 5140 52740 5196 52796
rect 5196 52740 5200 52796
rect 5136 52736 5200 52740
rect 5216 52796 5280 52800
rect 5216 52740 5220 52796
rect 5220 52740 5276 52796
rect 5276 52740 5280 52796
rect 5216 52736 5280 52740
rect 5296 52796 5360 52800
rect 5296 52740 5300 52796
rect 5300 52740 5356 52796
rect 5356 52740 5360 52796
rect 5296 52736 5360 52740
rect 5376 52796 5440 52800
rect 5376 52740 5380 52796
rect 5380 52740 5436 52796
rect 5436 52740 5440 52796
rect 5376 52736 5440 52740
rect 35856 52796 35920 52800
rect 35856 52740 35860 52796
rect 35860 52740 35916 52796
rect 35916 52740 35920 52796
rect 35856 52736 35920 52740
rect 35936 52796 36000 52800
rect 35936 52740 35940 52796
rect 35940 52740 35996 52796
rect 35996 52740 36000 52796
rect 35936 52736 36000 52740
rect 36016 52796 36080 52800
rect 36016 52740 36020 52796
rect 36020 52740 36076 52796
rect 36076 52740 36080 52796
rect 36016 52736 36080 52740
rect 36096 52796 36160 52800
rect 36096 52740 36100 52796
rect 36100 52740 36156 52796
rect 36156 52740 36160 52796
rect 36096 52736 36160 52740
rect 66576 52796 66640 52800
rect 66576 52740 66580 52796
rect 66580 52740 66636 52796
rect 66636 52740 66640 52796
rect 66576 52736 66640 52740
rect 66656 52796 66720 52800
rect 66656 52740 66660 52796
rect 66660 52740 66716 52796
rect 66716 52740 66720 52796
rect 66656 52736 66720 52740
rect 66736 52796 66800 52800
rect 66736 52740 66740 52796
rect 66740 52740 66796 52796
rect 66796 52740 66800 52796
rect 66736 52736 66800 52740
rect 66816 52796 66880 52800
rect 66816 52740 66820 52796
rect 66820 52740 66876 52796
rect 66876 52740 66880 52796
rect 66816 52736 66880 52740
rect 5796 52252 5860 52256
rect 5796 52196 5800 52252
rect 5800 52196 5856 52252
rect 5856 52196 5860 52252
rect 5796 52192 5860 52196
rect 5876 52252 5940 52256
rect 5876 52196 5880 52252
rect 5880 52196 5936 52252
rect 5936 52196 5940 52252
rect 5876 52192 5940 52196
rect 5956 52252 6020 52256
rect 5956 52196 5960 52252
rect 5960 52196 6016 52252
rect 6016 52196 6020 52252
rect 5956 52192 6020 52196
rect 6036 52252 6100 52256
rect 6036 52196 6040 52252
rect 6040 52196 6096 52252
rect 6096 52196 6100 52252
rect 6036 52192 6100 52196
rect 36516 52252 36580 52256
rect 36516 52196 36520 52252
rect 36520 52196 36576 52252
rect 36576 52196 36580 52252
rect 36516 52192 36580 52196
rect 36596 52252 36660 52256
rect 36596 52196 36600 52252
rect 36600 52196 36656 52252
rect 36656 52196 36660 52252
rect 36596 52192 36660 52196
rect 36676 52252 36740 52256
rect 36676 52196 36680 52252
rect 36680 52196 36736 52252
rect 36736 52196 36740 52252
rect 36676 52192 36740 52196
rect 36756 52252 36820 52256
rect 36756 52196 36760 52252
rect 36760 52196 36816 52252
rect 36816 52196 36820 52252
rect 36756 52192 36820 52196
rect 67236 52252 67300 52256
rect 67236 52196 67240 52252
rect 67240 52196 67296 52252
rect 67296 52196 67300 52252
rect 67236 52192 67300 52196
rect 67316 52252 67380 52256
rect 67316 52196 67320 52252
rect 67320 52196 67376 52252
rect 67376 52196 67380 52252
rect 67316 52192 67380 52196
rect 67396 52252 67460 52256
rect 67396 52196 67400 52252
rect 67400 52196 67456 52252
rect 67456 52196 67460 52252
rect 67396 52192 67460 52196
rect 67476 52252 67540 52256
rect 67476 52196 67480 52252
rect 67480 52196 67536 52252
rect 67536 52196 67540 52252
rect 67476 52192 67540 52196
rect 5136 51708 5200 51712
rect 5136 51652 5140 51708
rect 5140 51652 5196 51708
rect 5196 51652 5200 51708
rect 5136 51648 5200 51652
rect 5216 51708 5280 51712
rect 5216 51652 5220 51708
rect 5220 51652 5276 51708
rect 5276 51652 5280 51708
rect 5216 51648 5280 51652
rect 5296 51708 5360 51712
rect 5296 51652 5300 51708
rect 5300 51652 5356 51708
rect 5356 51652 5360 51708
rect 5296 51648 5360 51652
rect 5376 51708 5440 51712
rect 5376 51652 5380 51708
rect 5380 51652 5436 51708
rect 5436 51652 5440 51708
rect 5376 51648 5440 51652
rect 35856 51708 35920 51712
rect 35856 51652 35860 51708
rect 35860 51652 35916 51708
rect 35916 51652 35920 51708
rect 35856 51648 35920 51652
rect 35936 51708 36000 51712
rect 35936 51652 35940 51708
rect 35940 51652 35996 51708
rect 35996 51652 36000 51708
rect 35936 51648 36000 51652
rect 36016 51708 36080 51712
rect 36016 51652 36020 51708
rect 36020 51652 36076 51708
rect 36076 51652 36080 51708
rect 36016 51648 36080 51652
rect 36096 51708 36160 51712
rect 36096 51652 36100 51708
rect 36100 51652 36156 51708
rect 36156 51652 36160 51708
rect 36096 51648 36160 51652
rect 66576 51708 66640 51712
rect 66576 51652 66580 51708
rect 66580 51652 66636 51708
rect 66636 51652 66640 51708
rect 66576 51648 66640 51652
rect 66656 51708 66720 51712
rect 66656 51652 66660 51708
rect 66660 51652 66716 51708
rect 66716 51652 66720 51708
rect 66656 51648 66720 51652
rect 66736 51708 66800 51712
rect 66736 51652 66740 51708
rect 66740 51652 66796 51708
rect 66796 51652 66800 51708
rect 66736 51648 66800 51652
rect 66816 51708 66880 51712
rect 66816 51652 66820 51708
rect 66820 51652 66876 51708
rect 66876 51652 66880 51708
rect 66816 51648 66880 51652
rect 5796 51164 5860 51168
rect 5796 51108 5800 51164
rect 5800 51108 5856 51164
rect 5856 51108 5860 51164
rect 5796 51104 5860 51108
rect 5876 51164 5940 51168
rect 5876 51108 5880 51164
rect 5880 51108 5936 51164
rect 5936 51108 5940 51164
rect 5876 51104 5940 51108
rect 5956 51164 6020 51168
rect 5956 51108 5960 51164
rect 5960 51108 6016 51164
rect 6016 51108 6020 51164
rect 5956 51104 6020 51108
rect 6036 51164 6100 51168
rect 6036 51108 6040 51164
rect 6040 51108 6096 51164
rect 6096 51108 6100 51164
rect 6036 51104 6100 51108
rect 36516 51164 36580 51168
rect 36516 51108 36520 51164
rect 36520 51108 36576 51164
rect 36576 51108 36580 51164
rect 36516 51104 36580 51108
rect 36596 51164 36660 51168
rect 36596 51108 36600 51164
rect 36600 51108 36656 51164
rect 36656 51108 36660 51164
rect 36596 51104 36660 51108
rect 36676 51164 36740 51168
rect 36676 51108 36680 51164
rect 36680 51108 36736 51164
rect 36736 51108 36740 51164
rect 36676 51104 36740 51108
rect 36756 51164 36820 51168
rect 36756 51108 36760 51164
rect 36760 51108 36816 51164
rect 36816 51108 36820 51164
rect 36756 51104 36820 51108
rect 67236 51164 67300 51168
rect 67236 51108 67240 51164
rect 67240 51108 67296 51164
rect 67296 51108 67300 51164
rect 67236 51104 67300 51108
rect 67316 51164 67380 51168
rect 67316 51108 67320 51164
rect 67320 51108 67376 51164
rect 67376 51108 67380 51164
rect 67316 51104 67380 51108
rect 67396 51164 67460 51168
rect 67396 51108 67400 51164
rect 67400 51108 67456 51164
rect 67456 51108 67460 51164
rect 67396 51104 67460 51108
rect 67476 51164 67540 51168
rect 67476 51108 67480 51164
rect 67480 51108 67536 51164
rect 67536 51108 67540 51164
rect 67476 51104 67540 51108
rect 5136 50620 5200 50624
rect 5136 50564 5140 50620
rect 5140 50564 5196 50620
rect 5196 50564 5200 50620
rect 5136 50560 5200 50564
rect 5216 50620 5280 50624
rect 5216 50564 5220 50620
rect 5220 50564 5276 50620
rect 5276 50564 5280 50620
rect 5216 50560 5280 50564
rect 5296 50620 5360 50624
rect 5296 50564 5300 50620
rect 5300 50564 5356 50620
rect 5356 50564 5360 50620
rect 5296 50560 5360 50564
rect 5376 50620 5440 50624
rect 5376 50564 5380 50620
rect 5380 50564 5436 50620
rect 5436 50564 5440 50620
rect 5376 50560 5440 50564
rect 35856 50620 35920 50624
rect 35856 50564 35860 50620
rect 35860 50564 35916 50620
rect 35916 50564 35920 50620
rect 35856 50560 35920 50564
rect 35936 50620 36000 50624
rect 35936 50564 35940 50620
rect 35940 50564 35996 50620
rect 35996 50564 36000 50620
rect 35936 50560 36000 50564
rect 36016 50620 36080 50624
rect 36016 50564 36020 50620
rect 36020 50564 36076 50620
rect 36076 50564 36080 50620
rect 36016 50560 36080 50564
rect 36096 50620 36160 50624
rect 36096 50564 36100 50620
rect 36100 50564 36156 50620
rect 36156 50564 36160 50620
rect 36096 50560 36160 50564
rect 66576 50620 66640 50624
rect 66576 50564 66580 50620
rect 66580 50564 66636 50620
rect 66636 50564 66640 50620
rect 66576 50560 66640 50564
rect 66656 50620 66720 50624
rect 66656 50564 66660 50620
rect 66660 50564 66716 50620
rect 66716 50564 66720 50620
rect 66656 50560 66720 50564
rect 66736 50620 66800 50624
rect 66736 50564 66740 50620
rect 66740 50564 66796 50620
rect 66796 50564 66800 50620
rect 66736 50560 66800 50564
rect 66816 50620 66880 50624
rect 66816 50564 66820 50620
rect 66820 50564 66876 50620
rect 66876 50564 66880 50620
rect 66816 50560 66880 50564
rect 5796 50076 5860 50080
rect 5796 50020 5800 50076
rect 5800 50020 5856 50076
rect 5856 50020 5860 50076
rect 5796 50016 5860 50020
rect 5876 50076 5940 50080
rect 5876 50020 5880 50076
rect 5880 50020 5936 50076
rect 5936 50020 5940 50076
rect 5876 50016 5940 50020
rect 5956 50076 6020 50080
rect 5956 50020 5960 50076
rect 5960 50020 6016 50076
rect 6016 50020 6020 50076
rect 5956 50016 6020 50020
rect 6036 50076 6100 50080
rect 6036 50020 6040 50076
rect 6040 50020 6096 50076
rect 6096 50020 6100 50076
rect 6036 50016 6100 50020
rect 36516 50076 36580 50080
rect 36516 50020 36520 50076
rect 36520 50020 36576 50076
rect 36576 50020 36580 50076
rect 36516 50016 36580 50020
rect 36596 50076 36660 50080
rect 36596 50020 36600 50076
rect 36600 50020 36656 50076
rect 36656 50020 36660 50076
rect 36596 50016 36660 50020
rect 36676 50076 36740 50080
rect 36676 50020 36680 50076
rect 36680 50020 36736 50076
rect 36736 50020 36740 50076
rect 36676 50016 36740 50020
rect 36756 50076 36820 50080
rect 36756 50020 36760 50076
rect 36760 50020 36816 50076
rect 36816 50020 36820 50076
rect 36756 50016 36820 50020
rect 67236 50076 67300 50080
rect 67236 50020 67240 50076
rect 67240 50020 67296 50076
rect 67296 50020 67300 50076
rect 67236 50016 67300 50020
rect 67316 50076 67380 50080
rect 67316 50020 67320 50076
rect 67320 50020 67376 50076
rect 67376 50020 67380 50076
rect 67316 50016 67380 50020
rect 67396 50076 67460 50080
rect 67396 50020 67400 50076
rect 67400 50020 67456 50076
rect 67456 50020 67460 50076
rect 67396 50016 67460 50020
rect 67476 50076 67540 50080
rect 67476 50020 67480 50076
rect 67480 50020 67536 50076
rect 67536 50020 67540 50076
rect 67476 50016 67540 50020
rect 5136 49532 5200 49536
rect 5136 49476 5140 49532
rect 5140 49476 5196 49532
rect 5196 49476 5200 49532
rect 5136 49472 5200 49476
rect 5216 49532 5280 49536
rect 5216 49476 5220 49532
rect 5220 49476 5276 49532
rect 5276 49476 5280 49532
rect 5216 49472 5280 49476
rect 5296 49532 5360 49536
rect 5296 49476 5300 49532
rect 5300 49476 5356 49532
rect 5356 49476 5360 49532
rect 5296 49472 5360 49476
rect 5376 49532 5440 49536
rect 5376 49476 5380 49532
rect 5380 49476 5436 49532
rect 5436 49476 5440 49532
rect 5376 49472 5440 49476
rect 35856 49532 35920 49536
rect 35856 49476 35860 49532
rect 35860 49476 35916 49532
rect 35916 49476 35920 49532
rect 35856 49472 35920 49476
rect 35936 49532 36000 49536
rect 35936 49476 35940 49532
rect 35940 49476 35996 49532
rect 35996 49476 36000 49532
rect 35936 49472 36000 49476
rect 36016 49532 36080 49536
rect 36016 49476 36020 49532
rect 36020 49476 36076 49532
rect 36076 49476 36080 49532
rect 36016 49472 36080 49476
rect 36096 49532 36160 49536
rect 36096 49476 36100 49532
rect 36100 49476 36156 49532
rect 36156 49476 36160 49532
rect 36096 49472 36160 49476
rect 66576 49532 66640 49536
rect 66576 49476 66580 49532
rect 66580 49476 66636 49532
rect 66636 49476 66640 49532
rect 66576 49472 66640 49476
rect 66656 49532 66720 49536
rect 66656 49476 66660 49532
rect 66660 49476 66716 49532
rect 66716 49476 66720 49532
rect 66656 49472 66720 49476
rect 66736 49532 66800 49536
rect 66736 49476 66740 49532
rect 66740 49476 66796 49532
rect 66796 49476 66800 49532
rect 66736 49472 66800 49476
rect 66816 49532 66880 49536
rect 66816 49476 66820 49532
rect 66820 49476 66876 49532
rect 66876 49476 66880 49532
rect 66816 49472 66880 49476
rect 5796 48988 5860 48992
rect 5796 48932 5800 48988
rect 5800 48932 5856 48988
rect 5856 48932 5860 48988
rect 5796 48928 5860 48932
rect 5876 48988 5940 48992
rect 5876 48932 5880 48988
rect 5880 48932 5936 48988
rect 5936 48932 5940 48988
rect 5876 48928 5940 48932
rect 5956 48988 6020 48992
rect 5956 48932 5960 48988
rect 5960 48932 6016 48988
rect 6016 48932 6020 48988
rect 5956 48928 6020 48932
rect 6036 48988 6100 48992
rect 6036 48932 6040 48988
rect 6040 48932 6096 48988
rect 6096 48932 6100 48988
rect 6036 48928 6100 48932
rect 36516 48988 36580 48992
rect 36516 48932 36520 48988
rect 36520 48932 36576 48988
rect 36576 48932 36580 48988
rect 36516 48928 36580 48932
rect 36596 48988 36660 48992
rect 36596 48932 36600 48988
rect 36600 48932 36656 48988
rect 36656 48932 36660 48988
rect 36596 48928 36660 48932
rect 36676 48988 36740 48992
rect 36676 48932 36680 48988
rect 36680 48932 36736 48988
rect 36736 48932 36740 48988
rect 36676 48928 36740 48932
rect 36756 48988 36820 48992
rect 36756 48932 36760 48988
rect 36760 48932 36816 48988
rect 36816 48932 36820 48988
rect 36756 48928 36820 48932
rect 67236 48988 67300 48992
rect 67236 48932 67240 48988
rect 67240 48932 67296 48988
rect 67296 48932 67300 48988
rect 67236 48928 67300 48932
rect 67316 48988 67380 48992
rect 67316 48932 67320 48988
rect 67320 48932 67376 48988
rect 67376 48932 67380 48988
rect 67316 48928 67380 48932
rect 67396 48988 67460 48992
rect 67396 48932 67400 48988
rect 67400 48932 67456 48988
rect 67456 48932 67460 48988
rect 67396 48928 67460 48932
rect 67476 48988 67540 48992
rect 67476 48932 67480 48988
rect 67480 48932 67536 48988
rect 67536 48932 67540 48988
rect 67476 48928 67540 48932
rect 5136 48444 5200 48448
rect 5136 48388 5140 48444
rect 5140 48388 5196 48444
rect 5196 48388 5200 48444
rect 5136 48384 5200 48388
rect 5216 48444 5280 48448
rect 5216 48388 5220 48444
rect 5220 48388 5276 48444
rect 5276 48388 5280 48444
rect 5216 48384 5280 48388
rect 5296 48444 5360 48448
rect 5296 48388 5300 48444
rect 5300 48388 5356 48444
rect 5356 48388 5360 48444
rect 5296 48384 5360 48388
rect 5376 48444 5440 48448
rect 5376 48388 5380 48444
rect 5380 48388 5436 48444
rect 5436 48388 5440 48444
rect 5376 48384 5440 48388
rect 35856 48444 35920 48448
rect 35856 48388 35860 48444
rect 35860 48388 35916 48444
rect 35916 48388 35920 48444
rect 35856 48384 35920 48388
rect 35936 48444 36000 48448
rect 35936 48388 35940 48444
rect 35940 48388 35996 48444
rect 35996 48388 36000 48444
rect 35936 48384 36000 48388
rect 36016 48444 36080 48448
rect 36016 48388 36020 48444
rect 36020 48388 36076 48444
rect 36076 48388 36080 48444
rect 36016 48384 36080 48388
rect 36096 48444 36160 48448
rect 36096 48388 36100 48444
rect 36100 48388 36156 48444
rect 36156 48388 36160 48444
rect 36096 48384 36160 48388
rect 66576 48444 66640 48448
rect 66576 48388 66580 48444
rect 66580 48388 66636 48444
rect 66636 48388 66640 48444
rect 66576 48384 66640 48388
rect 66656 48444 66720 48448
rect 66656 48388 66660 48444
rect 66660 48388 66716 48444
rect 66716 48388 66720 48444
rect 66656 48384 66720 48388
rect 66736 48444 66800 48448
rect 66736 48388 66740 48444
rect 66740 48388 66796 48444
rect 66796 48388 66800 48444
rect 66736 48384 66800 48388
rect 66816 48444 66880 48448
rect 66816 48388 66820 48444
rect 66820 48388 66876 48444
rect 66876 48388 66880 48444
rect 66816 48384 66880 48388
rect 5796 47900 5860 47904
rect 5796 47844 5800 47900
rect 5800 47844 5856 47900
rect 5856 47844 5860 47900
rect 5796 47840 5860 47844
rect 5876 47900 5940 47904
rect 5876 47844 5880 47900
rect 5880 47844 5936 47900
rect 5936 47844 5940 47900
rect 5876 47840 5940 47844
rect 5956 47900 6020 47904
rect 5956 47844 5960 47900
rect 5960 47844 6016 47900
rect 6016 47844 6020 47900
rect 5956 47840 6020 47844
rect 6036 47900 6100 47904
rect 6036 47844 6040 47900
rect 6040 47844 6096 47900
rect 6096 47844 6100 47900
rect 6036 47840 6100 47844
rect 36516 47900 36580 47904
rect 36516 47844 36520 47900
rect 36520 47844 36576 47900
rect 36576 47844 36580 47900
rect 36516 47840 36580 47844
rect 36596 47900 36660 47904
rect 36596 47844 36600 47900
rect 36600 47844 36656 47900
rect 36656 47844 36660 47900
rect 36596 47840 36660 47844
rect 36676 47900 36740 47904
rect 36676 47844 36680 47900
rect 36680 47844 36736 47900
rect 36736 47844 36740 47900
rect 36676 47840 36740 47844
rect 36756 47900 36820 47904
rect 36756 47844 36760 47900
rect 36760 47844 36816 47900
rect 36816 47844 36820 47900
rect 36756 47840 36820 47844
rect 67236 47900 67300 47904
rect 67236 47844 67240 47900
rect 67240 47844 67296 47900
rect 67296 47844 67300 47900
rect 67236 47840 67300 47844
rect 67316 47900 67380 47904
rect 67316 47844 67320 47900
rect 67320 47844 67376 47900
rect 67376 47844 67380 47900
rect 67316 47840 67380 47844
rect 67396 47900 67460 47904
rect 67396 47844 67400 47900
rect 67400 47844 67456 47900
rect 67456 47844 67460 47900
rect 67396 47840 67460 47844
rect 67476 47900 67540 47904
rect 67476 47844 67480 47900
rect 67480 47844 67536 47900
rect 67536 47844 67540 47900
rect 67476 47840 67540 47844
rect 5136 47356 5200 47360
rect 5136 47300 5140 47356
rect 5140 47300 5196 47356
rect 5196 47300 5200 47356
rect 5136 47296 5200 47300
rect 5216 47356 5280 47360
rect 5216 47300 5220 47356
rect 5220 47300 5276 47356
rect 5276 47300 5280 47356
rect 5216 47296 5280 47300
rect 5296 47356 5360 47360
rect 5296 47300 5300 47356
rect 5300 47300 5356 47356
rect 5356 47300 5360 47356
rect 5296 47296 5360 47300
rect 5376 47356 5440 47360
rect 5376 47300 5380 47356
rect 5380 47300 5436 47356
rect 5436 47300 5440 47356
rect 5376 47296 5440 47300
rect 35856 47356 35920 47360
rect 35856 47300 35860 47356
rect 35860 47300 35916 47356
rect 35916 47300 35920 47356
rect 35856 47296 35920 47300
rect 35936 47356 36000 47360
rect 35936 47300 35940 47356
rect 35940 47300 35996 47356
rect 35996 47300 36000 47356
rect 35936 47296 36000 47300
rect 36016 47356 36080 47360
rect 36016 47300 36020 47356
rect 36020 47300 36076 47356
rect 36076 47300 36080 47356
rect 36016 47296 36080 47300
rect 36096 47356 36160 47360
rect 36096 47300 36100 47356
rect 36100 47300 36156 47356
rect 36156 47300 36160 47356
rect 36096 47296 36160 47300
rect 66576 47356 66640 47360
rect 66576 47300 66580 47356
rect 66580 47300 66636 47356
rect 66636 47300 66640 47356
rect 66576 47296 66640 47300
rect 66656 47356 66720 47360
rect 66656 47300 66660 47356
rect 66660 47300 66716 47356
rect 66716 47300 66720 47356
rect 66656 47296 66720 47300
rect 66736 47356 66800 47360
rect 66736 47300 66740 47356
rect 66740 47300 66796 47356
rect 66796 47300 66800 47356
rect 66736 47296 66800 47300
rect 66816 47356 66880 47360
rect 66816 47300 66820 47356
rect 66820 47300 66876 47356
rect 66876 47300 66880 47356
rect 66816 47296 66880 47300
rect 5796 46812 5860 46816
rect 5796 46756 5800 46812
rect 5800 46756 5856 46812
rect 5856 46756 5860 46812
rect 5796 46752 5860 46756
rect 5876 46812 5940 46816
rect 5876 46756 5880 46812
rect 5880 46756 5936 46812
rect 5936 46756 5940 46812
rect 5876 46752 5940 46756
rect 5956 46812 6020 46816
rect 5956 46756 5960 46812
rect 5960 46756 6016 46812
rect 6016 46756 6020 46812
rect 5956 46752 6020 46756
rect 6036 46812 6100 46816
rect 6036 46756 6040 46812
rect 6040 46756 6096 46812
rect 6096 46756 6100 46812
rect 6036 46752 6100 46756
rect 36516 46812 36580 46816
rect 36516 46756 36520 46812
rect 36520 46756 36576 46812
rect 36576 46756 36580 46812
rect 36516 46752 36580 46756
rect 36596 46812 36660 46816
rect 36596 46756 36600 46812
rect 36600 46756 36656 46812
rect 36656 46756 36660 46812
rect 36596 46752 36660 46756
rect 36676 46812 36740 46816
rect 36676 46756 36680 46812
rect 36680 46756 36736 46812
rect 36736 46756 36740 46812
rect 36676 46752 36740 46756
rect 36756 46812 36820 46816
rect 36756 46756 36760 46812
rect 36760 46756 36816 46812
rect 36816 46756 36820 46812
rect 36756 46752 36820 46756
rect 67236 46812 67300 46816
rect 67236 46756 67240 46812
rect 67240 46756 67296 46812
rect 67296 46756 67300 46812
rect 67236 46752 67300 46756
rect 67316 46812 67380 46816
rect 67316 46756 67320 46812
rect 67320 46756 67376 46812
rect 67376 46756 67380 46812
rect 67316 46752 67380 46756
rect 67396 46812 67460 46816
rect 67396 46756 67400 46812
rect 67400 46756 67456 46812
rect 67456 46756 67460 46812
rect 67396 46752 67460 46756
rect 67476 46812 67540 46816
rect 67476 46756 67480 46812
rect 67480 46756 67536 46812
rect 67536 46756 67540 46812
rect 67476 46752 67540 46756
rect 5136 46268 5200 46272
rect 5136 46212 5140 46268
rect 5140 46212 5196 46268
rect 5196 46212 5200 46268
rect 5136 46208 5200 46212
rect 5216 46268 5280 46272
rect 5216 46212 5220 46268
rect 5220 46212 5276 46268
rect 5276 46212 5280 46268
rect 5216 46208 5280 46212
rect 5296 46268 5360 46272
rect 5296 46212 5300 46268
rect 5300 46212 5356 46268
rect 5356 46212 5360 46268
rect 5296 46208 5360 46212
rect 5376 46268 5440 46272
rect 5376 46212 5380 46268
rect 5380 46212 5436 46268
rect 5436 46212 5440 46268
rect 5376 46208 5440 46212
rect 35856 46268 35920 46272
rect 35856 46212 35860 46268
rect 35860 46212 35916 46268
rect 35916 46212 35920 46268
rect 35856 46208 35920 46212
rect 35936 46268 36000 46272
rect 35936 46212 35940 46268
rect 35940 46212 35996 46268
rect 35996 46212 36000 46268
rect 35936 46208 36000 46212
rect 36016 46268 36080 46272
rect 36016 46212 36020 46268
rect 36020 46212 36076 46268
rect 36076 46212 36080 46268
rect 36016 46208 36080 46212
rect 36096 46268 36160 46272
rect 36096 46212 36100 46268
rect 36100 46212 36156 46268
rect 36156 46212 36160 46268
rect 36096 46208 36160 46212
rect 66576 46268 66640 46272
rect 66576 46212 66580 46268
rect 66580 46212 66636 46268
rect 66636 46212 66640 46268
rect 66576 46208 66640 46212
rect 66656 46268 66720 46272
rect 66656 46212 66660 46268
rect 66660 46212 66716 46268
rect 66716 46212 66720 46268
rect 66656 46208 66720 46212
rect 66736 46268 66800 46272
rect 66736 46212 66740 46268
rect 66740 46212 66796 46268
rect 66796 46212 66800 46268
rect 66736 46208 66800 46212
rect 66816 46268 66880 46272
rect 66816 46212 66820 46268
rect 66820 46212 66876 46268
rect 66876 46212 66880 46268
rect 66816 46208 66880 46212
rect 5796 45724 5860 45728
rect 5796 45668 5800 45724
rect 5800 45668 5856 45724
rect 5856 45668 5860 45724
rect 5796 45664 5860 45668
rect 5876 45724 5940 45728
rect 5876 45668 5880 45724
rect 5880 45668 5936 45724
rect 5936 45668 5940 45724
rect 5876 45664 5940 45668
rect 5956 45724 6020 45728
rect 5956 45668 5960 45724
rect 5960 45668 6016 45724
rect 6016 45668 6020 45724
rect 5956 45664 6020 45668
rect 6036 45724 6100 45728
rect 6036 45668 6040 45724
rect 6040 45668 6096 45724
rect 6096 45668 6100 45724
rect 6036 45664 6100 45668
rect 36516 45724 36580 45728
rect 36516 45668 36520 45724
rect 36520 45668 36576 45724
rect 36576 45668 36580 45724
rect 36516 45664 36580 45668
rect 36596 45724 36660 45728
rect 36596 45668 36600 45724
rect 36600 45668 36656 45724
rect 36656 45668 36660 45724
rect 36596 45664 36660 45668
rect 36676 45724 36740 45728
rect 36676 45668 36680 45724
rect 36680 45668 36736 45724
rect 36736 45668 36740 45724
rect 36676 45664 36740 45668
rect 36756 45724 36820 45728
rect 36756 45668 36760 45724
rect 36760 45668 36816 45724
rect 36816 45668 36820 45724
rect 36756 45664 36820 45668
rect 67236 45724 67300 45728
rect 67236 45668 67240 45724
rect 67240 45668 67296 45724
rect 67296 45668 67300 45724
rect 67236 45664 67300 45668
rect 67316 45724 67380 45728
rect 67316 45668 67320 45724
rect 67320 45668 67376 45724
rect 67376 45668 67380 45724
rect 67316 45664 67380 45668
rect 67396 45724 67460 45728
rect 67396 45668 67400 45724
rect 67400 45668 67456 45724
rect 67456 45668 67460 45724
rect 67396 45664 67460 45668
rect 67476 45724 67540 45728
rect 67476 45668 67480 45724
rect 67480 45668 67536 45724
rect 67536 45668 67540 45724
rect 67476 45664 67540 45668
rect 5136 45180 5200 45184
rect 5136 45124 5140 45180
rect 5140 45124 5196 45180
rect 5196 45124 5200 45180
rect 5136 45120 5200 45124
rect 5216 45180 5280 45184
rect 5216 45124 5220 45180
rect 5220 45124 5276 45180
rect 5276 45124 5280 45180
rect 5216 45120 5280 45124
rect 5296 45180 5360 45184
rect 5296 45124 5300 45180
rect 5300 45124 5356 45180
rect 5356 45124 5360 45180
rect 5296 45120 5360 45124
rect 5376 45180 5440 45184
rect 5376 45124 5380 45180
rect 5380 45124 5436 45180
rect 5436 45124 5440 45180
rect 5376 45120 5440 45124
rect 35856 45180 35920 45184
rect 35856 45124 35860 45180
rect 35860 45124 35916 45180
rect 35916 45124 35920 45180
rect 35856 45120 35920 45124
rect 35936 45180 36000 45184
rect 35936 45124 35940 45180
rect 35940 45124 35996 45180
rect 35996 45124 36000 45180
rect 35936 45120 36000 45124
rect 36016 45180 36080 45184
rect 36016 45124 36020 45180
rect 36020 45124 36076 45180
rect 36076 45124 36080 45180
rect 36016 45120 36080 45124
rect 36096 45180 36160 45184
rect 36096 45124 36100 45180
rect 36100 45124 36156 45180
rect 36156 45124 36160 45180
rect 36096 45120 36160 45124
rect 66576 45180 66640 45184
rect 66576 45124 66580 45180
rect 66580 45124 66636 45180
rect 66636 45124 66640 45180
rect 66576 45120 66640 45124
rect 66656 45180 66720 45184
rect 66656 45124 66660 45180
rect 66660 45124 66716 45180
rect 66716 45124 66720 45180
rect 66656 45120 66720 45124
rect 66736 45180 66800 45184
rect 66736 45124 66740 45180
rect 66740 45124 66796 45180
rect 66796 45124 66800 45180
rect 66736 45120 66800 45124
rect 66816 45180 66880 45184
rect 66816 45124 66820 45180
rect 66820 45124 66876 45180
rect 66876 45124 66880 45180
rect 66816 45120 66880 45124
rect 5796 44636 5860 44640
rect 5796 44580 5800 44636
rect 5800 44580 5856 44636
rect 5856 44580 5860 44636
rect 5796 44576 5860 44580
rect 5876 44636 5940 44640
rect 5876 44580 5880 44636
rect 5880 44580 5936 44636
rect 5936 44580 5940 44636
rect 5876 44576 5940 44580
rect 5956 44636 6020 44640
rect 5956 44580 5960 44636
rect 5960 44580 6016 44636
rect 6016 44580 6020 44636
rect 5956 44576 6020 44580
rect 6036 44636 6100 44640
rect 6036 44580 6040 44636
rect 6040 44580 6096 44636
rect 6096 44580 6100 44636
rect 6036 44576 6100 44580
rect 36516 44636 36580 44640
rect 36516 44580 36520 44636
rect 36520 44580 36576 44636
rect 36576 44580 36580 44636
rect 36516 44576 36580 44580
rect 36596 44636 36660 44640
rect 36596 44580 36600 44636
rect 36600 44580 36656 44636
rect 36656 44580 36660 44636
rect 36596 44576 36660 44580
rect 36676 44636 36740 44640
rect 36676 44580 36680 44636
rect 36680 44580 36736 44636
rect 36736 44580 36740 44636
rect 36676 44576 36740 44580
rect 36756 44636 36820 44640
rect 36756 44580 36760 44636
rect 36760 44580 36816 44636
rect 36816 44580 36820 44636
rect 36756 44576 36820 44580
rect 67236 44636 67300 44640
rect 67236 44580 67240 44636
rect 67240 44580 67296 44636
rect 67296 44580 67300 44636
rect 67236 44576 67300 44580
rect 67316 44636 67380 44640
rect 67316 44580 67320 44636
rect 67320 44580 67376 44636
rect 67376 44580 67380 44636
rect 67316 44576 67380 44580
rect 67396 44636 67460 44640
rect 67396 44580 67400 44636
rect 67400 44580 67456 44636
rect 67456 44580 67460 44636
rect 67396 44576 67460 44580
rect 67476 44636 67540 44640
rect 67476 44580 67480 44636
rect 67480 44580 67536 44636
rect 67536 44580 67540 44636
rect 67476 44576 67540 44580
rect 5136 44092 5200 44096
rect 5136 44036 5140 44092
rect 5140 44036 5196 44092
rect 5196 44036 5200 44092
rect 5136 44032 5200 44036
rect 5216 44092 5280 44096
rect 5216 44036 5220 44092
rect 5220 44036 5276 44092
rect 5276 44036 5280 44092
rect 5216 44032 5280 44036
rect 5296 44092 5360 44096
rect 5296 44036 5300 44092
rect 5300 44036 5356 44092
rect 5356 44036 5360 44092
rect 5296 44032 5360 44036
rect 5376 44092 5440 44096
rect 5376 44036 5380 44092
rect 5380 44036 5436 44092
rect 5436 44036 5440 44092
rect 5376 44032 5440 44036
rect 35856 44092 35920 44096
rect 35856 44036 35860 44092
rect 35860 44036 35916 44092
rect 35916 44036 35920 44092
rect 35856 44032 35920 44036
rect 35936 44092 36000 44096
rect 35936 44036 35940 44092
rect 35940 44036 35996 44092
rect 35996 44036 36000 44092
rect 35936 44032 36000 44036
rect 36016 44092 36080 44096
rect 36016 44036 36020 44092
rect 36020 44036 36076 44092
rect 36076 44036 36080 44092
rect 36016 44032 36080 44036
rect 36096 44092 36160 44096
rect 36096 44036 36100 44092
rect 36100 44036 36156 44092
rect 36156 44036 36160 44092
rect 36096 44032 36160 44036
rect 66576 44092 66640 44096
rect 66576 44036 66580 44092
rect 66580 44036 66636 44092
rect 66636 44036 66640 44092
rect 66576 44032 66640 44036
rect 66656 44092 66720 44096
rect 66656 44036 66660 44092
rect 66660 44036 66716 44092
rect 66716 44036 66720 44092
rect 66656 44032 66720 44036
rect 66736 44092 66800 44096
rect 66736 44036 66740 44092
rect 66740 44036 66796 44092
rect 66796 44036 66800 44092
rect 66736 44032 66800 44036
rect 66816 44092 66880 44096
rect 66816 44036 66820 44092
rect 66820 44036 66876 44092
rect 66876 44036 66880 44092
rect 66816 44032 66880 44036
rect 5796 43548 5860 43552
rect 5796 43492 5800 43548
rect 5800 43492 5856 43548
rect 5856 43492 5860 43548
rect 5796 43488 5860 43492
rect 5876 43548 5940 43552
rect 5876 43492 5880 43548
rect 5880 43492 5936 43548
rect 5936 43492 5940 43548
rect 5876 43488 5940 43492
rect 5956 43548 6020 43552
rect 5956 43492 5960 43548
rect 5960 43492 6016 43548
rect 6016 43492 6020 43548
rect 5956 43488 6020 43492
rect 6036 43548 6100 43552
rect 6036 43492 6040 43548
rect 6040 43492 6096 43548
rect 6096 43492 6100 43548
rect 6036 43488 6100 43492
rect 36516 43548 36580 43552
rect 36516 43492 36520 43548
rect 36520 43492 36576 43548
rect 36576 43492 36580 43548
rect 36516 43488 36580 43492
rect 36596 43548 36660 43552
rect 36596 43492 36600 43548
rect 36600 43492 36656 43548
rect 36656 43492 36660 43548
rect 36596 43488 36660 43492
rect 36676 43548 36740 43552
rect 36676 43492 36680 43548
rect 36680 43492 36736 43548
rect 36736 43492 36740 43548
rect 36676 43488 36740 43492
rect 36756 43548 36820 43552
rect 36756 43492 36760 43548
rect 36760 43492 36816 43548
rect 36816 43492 36820 43548
rect 36756 43488 36820 43492
rect 67236 43548 67300 43552
rect 67236 43492 67240 43548
rect 67240 43492 67296 43548
rect 67296 43492 67300 43548
rect 67236 43488 67300 43492
rect 67316 43548 67380 43552
rect 67316 43492 67320 43548
rect 67320 43492 67376 43548
rect 67376 43492 67380 43548
rect 67316 43488 67380 43492
rect 67396 43548 67460 43552
rect 67396 43492 67400 43548
rect 67400 43492 67456 43548
rect 67456 43492 67460 43548
rect 67396 43488 67460 43492
rect 67476 43548 67540 43552
rect 67476 43492 67480 43548
rect 67480 43492 67536 43548
rect 67536 43492 67540 43548
rect 67476 43488 67540 43492
rect 5136 43004 5200 43008
rect 5136 42948 5140 43004
rect 5140 42948 5196 43004
rect 5196 42948 5200 43004
rect 5136 42944 5200 42948
rect 5216 43004 5280 43008
rect 5216 42948 5220 43004
rect 5220 42948 5276 43004
rect 5276 42948 5280 43004
rect 5216 42944 5280 42948
rect 5296 43004 5360 43008
rect 5296 42948 5300 43004
rect 5300 42948 5356 43004
rect 5356 42948 5360 43004
rect 5296 42944 5360 42948
rect 5376 43004 5440 43008
rect 5376 42948 5380 43004
rect 5380 42948 5436 43004
rect 5436 42948 5440 43004
rect 5376 42944 5440 42948
rect 35856 43004 35920 43008
rect 35856 42948 35860 43004
rect 35860 42948 35916 43004
rect 35916 42948 35920 43004
rect 35856 42944 35920 42948
rect 35936 43004 36000 43008
rect 35936 42948 35940 43004
rect 35940 42948 35996 43004
rect 35996 42948 36000 43004
rect 35936 42944 36000 42948
rect 36016 43004 36080 43008
rect 36016 42948 36020 43004
rect 36020 42948 36076 43004
rect 36076 42948 36080 43004
rect 36016 42944 36080 42948
rect 36096 43004 36160 43008
rect 36096 42948 36100 43004
rect 36100 42948 36156 43004
rect 36156 42948 36160 43004
rect 36096 42944 36160 42948
rect 66576 43004 66640 43008
rect 66576 42948 66580 43004
rect 66580 42948 66636 43004
rect 66636 42948 66640 43004
rect 66576 42944 66640 42948
rect 66656 43004 66720 43008
rect 66656 42948 66660 43004
rect 66660 42948 66716 43004
rect 66716 42948 66720 43004
rect 66656 42944 66720 42948
rect 66736 43004 66800 43008
rect 66736 42948 66740 43004
rect 66740 42948 66796 43004
rect 66796 42948 66800 43004
rect 66736 42944 66800 42948
rect 66816 43004 66880 43008
rect 66816 42948 66820 43004
rect 66820 42948 66876 43004
rect 66876 42948 66880 43004
rect 66816 42944 66880 42948
rect 5796 42460 5860 42464
rect 5796 42404 5800 42460
rect 5800 42404 5856 42460
rect 5856 42404 5860 42460
rect 5796 42400 5860 42404
rect 5876 42460 5940 42464
rect 5876 42404 5880 42460
rect 5880 42404 5936 42460
rect 5936 42404 5940 42460
rect 5876 42400 5940 42404
rect 5956 42460 6020 42464
rect 5956 42404 5960 42460
rect 5960 42404 6016 42460
rect 6016 42404 6020 42460
rect 5956 42400 6020 42404
rect 6036 42460 6100 42464
rect 6036 42404 6040 42460
rect 6040 42404 6096 42460
rect 6096 42404 6100 42460
rect 6036 42400 6100 42404
rect 36516 42460 36580 42464
rect 36516 42404 36520 42460
rect 36520 42404 36576 42460
rect 36576 42404 36580 42460
rect 36516 42400 36580 42404
rect 36596 42460 36660 42464
rect 36596 42404 36600 42460
rect 36600 42404 36656 42460
rect 36656 42404 36660 42460
rect 36596 42400 36660 42404
rect 36676 42460 36740 42464
rect 36676 42404 36680 42460
rect 36680 42404 36736 42460
rect 36736 42404 36740 42460
rect 36676 42400 36740 42404
rect 36756 42460 36820 42464
rect 36756 42404 36760 42460
rect 36760 42404 36816 42460
rect 36816 42404 36820 42460
rect 36756 42400 36820 42404
rect 67236 42460 67300 42464
rect 67236 42404 67240 42460
rect 67240 42404 67296 42460
rect 67296 42404 67300 42460
rect 67236 42400 67300 42404
rect 67316 42460 67380 42464
rect 67316 42404 67320 42460
rect 67320 42404 67376 42460
rect 67376 42404 67380 42460
rect 67316 42400 67380 42404
rect 67396 42460 67460 42464
rect 67396 42404 67400 42460
rect 67400 42404 67456 42460
rect 67456 42404 67460 42460
rect 67396 42400 67460 42404
rect 67476 42460 67540 42464
rect 67476 42404 67480 42460
rect 67480 42404 67536 42460
rect 67536 42404 67540 42460
rect 67476 42400 67540 42404
rect 5136 41916 5200 41920
rect 5136 41860 5140 41916
rect 5140 41860 5196 41916
rect 5196 41860 5200 41916
rect 5136 41856 5200 41860
rect 5216 41916 5280 41920
rect 5216 41860 5220 41916
rect 5220 41860 5276 41916
rect 5276 41860 5280 41916
rect 5216 41856 5280 41860
rect 5296 41916 5360 41920
rect 5296 41860 5300 41916
rect 5300 41860 5356 41916
rect 5356 41860 5360 41916
rect 5296 41856 5360 41860
rect 5376 41916 5440 41920
rect 5376 41860 5380 41916
rect 5380 41860 5436 41916
rect 5436 41860 5440 41916
rect 5376 41856 5440 41860
rect 35856 41916 35920 41920
rect 35856 41860 35860 41916
rect 35860 41860 35916 41916
rect 35916 41860 35920 41916
rect 35856 41856 35920 41860
rect 35936 41916 36000 41920
rect 35936 41860 35940 41916
rect 35940 41860 35996 41916
rect 35996 41860 36000 41916
rect 35936 41856 36000 41860
rect 36016 41916 36080 41920
rect 36016 41860 36020 41916
rect 36020 41860 36076 41916
rect 36076 41860 36080 41916
rect 36016 41856 36080 41860
rect 36096 41916 36160 41920
rect 36096 41860 36100 41916
rect 36100 41860 36156 41916
rect 36156 41860 36160 41916
rect 36096 41856 36160 41860
rect 66576 41916 66640 41920
rect 66576 41860 66580 41916
rect 66580 41860 66636 41916
rect 66636 41860 66640 41916
rect 66576 41856 66640 41860
rect 66656 41916 66720 41920
rect 66656 41860 66660 41916
rect 66660 41860 66716 41916
rect 66716 41860 66720 41916
rect 66656 41856 66720 41860
rect 66736 41916 66800 41920
rect 66736 41860 66740 41916
rect 66740 41860 66796 41916
rect 66796 41860 66800 41916
rect 66736 41856 66800 41860
rect 66816 41916 66880 41920
rect 66816 41860 66820 41916
rect 66820 41860 66876 41916
rect 66876 41860 66880 41916
rect 66816 41856 66880 41860
rect 5796 41372 5860 41376
rect 5796 41316 5800 41372
rect 5800 41316 5856 41372
rect 5856 41316 5860 41372
rect 5796 41312 5860 41316
rect 5876 41372 5940 41376
rect 5876 41316 5880 41372
rect 5880 41316 5936 41372
rect 5936 41316 5940 41372
rect 5876 41312 5940 41316
rect 5956 41372 6020 41376
rect 5956 41316 5960 41372
rect 5960 41316 6016 41372
rect 6016 41316 6020 41372
rect 5956 41312 6020 41316
rect 6036 41372 6100 41376
rect 6036 41316 6040 41372
rect 6040 41316 6096 41372
rect 6096 41316 6100 41372
rect 6036 41312 6100 41316
rect 36516 41372 36580 41376
rect 36516 41316 36520 41372
rect 36520 41316 36576 41372
rect 36576 41316 36580 41372
rect 36516 41312 36580 41316
rect 36596 41372 36660 41376
rect 36596 41316 36600 41372
rect 36600 41316 36656 41372
rect 36656 41316 36660 41372
rect 36596 41312 36660 41316
rect 36676 41372 36740 41376
rect 36676 41316 36680 41372
rect 36680 41316 36736 41372
rect 36736 41316 36740 41372
rect 36676 41312 36740 41316
rect 36756 41372 36820 41376
rect 36756 41316 36760 41372
rect 36760 41316 36816 41372
rect 36816 41316 36820 41372
rect 36756 41312 36820 41316
rect 67236 41372 67300 41376
rect 67236 41316 67240 41372
rect 67240 41316 67296 41372
rect 67296 41316 67300 41372
rect 67236 41312 67300 41316
rect 67316 41372 67380 41376
rect 67316 41316 67320 41372
rect 67320 41316 67376 41372
rect 67376 41316 67380 41372
rect 67316 41312 67380 41316
rect 67396 41372 67460 41376
rect 67396 41316 67400 41372
rect 67400 41316 67456 41372
rect 67456 41316 67460 41372
rect 67396 41312 67460 41316
rect 67476 41372 67540 41376
rect 67476 41316 67480 41372
rect 67480 41316 67536 41372
rect 67536 41316 67540 41372
rect 67476 41312 67540 41316
rect 5136 40828 5200 40832
rect 5136 40772 5140 40828
rect 5140 40772 5196 40828
rect 5196 40772 5200 40828
rect 5136 40768 5200 40772
rect 5216 40828 5280 40832
rect 5216 40772 5220 40828
rect 5220 40772 5276 40828
rect 5276 40772 5280 40828
rect 5216 40768 5280 40772
rect 5296 40828 5360 40832
rect 5296 40772 5300 40828
rect 5300 40772 5356 40828
rect 5356 40772 5360 40828
rect 5296 40768 5360 40772
rect 5376 40828 5440 40832
rect 5376 40772 5380 40828
rect 5380 40772 5436 40828
rect 5436 40772 5440 40828
rect 5376 40768 5440 40772
rect 35856 40828 35920 40832
rect 35856 40772 35860 40828
rect 35860 40772 35916 40828
rect 35916 40772 35920 40828
rect 35856 40768 35920 40772
rect 35936 40828 36000 40832
rect 35936 40772 35940 40828
rect 35940 40772 35996 40828
rect 35996 40772 36000 40828
rect 35936 40768 36000 40772
rect 36016 40828 36080 40832
rect 36016 40772 36020 40828
rect 36020 40772 36076 40828
rect 36076 40772 36080 40828
rect 36016 40768 36080 40772
rect 36096 40828 36160 40832
rect 36096 40772 36100 40828
rect 36100 40772 36156 40828
rect 36156 40772 36160 40828
rect 36096 40768 36160 40772
rect 66576 40828 66640 40832
rect 66576 40772 66580 40828
rect 66580 40772 66636 40828
rect 66636 40772 66640 40828
rect 66576 40768 66640 40772
rect 66656 40828 66720 40832
rect 66656 40772 66660 40828
rect 66660 40772 66716 40828
rect 66716 40772 66720 40828
rect 66656 40768 66720 40772
rect 66736 40828 66800 40832
rect 66736 40772 66740 40828
rect 66740 40772 66796 40828
rect 66796 40772 66800 40828
rect 66736 40768 66800 40772
rect 66816 40828 66880 40832
rect 66816 40772 66820 40828
rect 66820 40772 66876 40828
rect 66876 40772 66880 40828
rect 66816 40768 66880 40772
rect 5796 40284 5860 40288
rect 5796 40228 5800 40284
rect 5800 40228 5856 40284
rect 5856 40228 5860 40284
rect 5796 40224 5860 40228
rect 5876 40284 5940 40288
rect 5876 40228 5880 40284
rect 5880 40228 5936 40284
rect 5936 40228 5940 40284
rect 5876 40224 5940 40228
rect 5956 40284 6020 40288
rect 5956 40228 5960 40284
rect 5960 40228 6016 40284
rect 6016 40228 6020 40284
rect 5956 40224 6020 40228
rect 6036 40284 6100 40288
rect 6036 40228 6040 40284
rect 6040 40228 6096 40284
rect 6096 40228 6100 40284
rect 6036 40224 6100 40228
rect 36516 40284 36580 40288
rect 36516 40228 36520 40284
rect 36520 40228 36576 40284
rect 36576 40228 36580 40284
rect 36516 40224 36580 40228
rect 36596 40284 36660 40288
rect 36596 40228 36600 40284
rect 36600 40228 36656 40284
rect 36656 40228 36660 40284
rect 36596 40224 36660 40228
rect 36676 40284 36740 40288
rect 36676 40228 36680 40284
rect 36680 40228 36736 40284
rect 36736 40228 36740 40284
rect 36676 40224 36740 40228
rect 36756 40284 36820 40288
rect 36756 40228 36760 40284
rect 36760 40228 36816 40284
rect 36816 40228 36820 40284
rect 36756 40224 36820 40228
rect 67236 40284 67300 40288
rect 67236 40228 67240 40284
rect 67240 40228 67296 40284
rect 67296 40228 67300 40284
rect 67236 40224 67300 40228
rect 67316 40284 67380 40288
rect 67316 40228 67320 40284
rect 67320 40228 67376 40284
rect 67376 40228 67380 40284
rect 67316 40224 67380 40228
rect 67396 40284 67460 40288
rect 67396 40228 67400 40284
rect 67400 40228 67456 40284
rect 67456 40228 67460 40284
rect 67396 40224 67460 40228
rect 67476 40284 67540 40288
rect 67476 40228 67480 40284
rect 67480 40228 67536 40284
rect 67536 40228 67540 40284
rect 67476 40224 67540 40228
rect 5136 39740 5200 39744
rect 5136 39684 5140 39740
rect 5140 39684 5196 39740
rect 5196 39684 5200 39740
rect 5136 39680 5200 39684
rect 5216 39740 5280 39744
rect 5216 39684 5220 39740
rect 5220 39684 5276 39740
rect 5276 39684 5280 39740
rect 5216 39680 5280 39684
rect 5296 39740 5360 39744
rect 5296 39684 5300 39740
rect 5300 39684 5356 39740
rect 5356 39684 5360 39740
rect 5296 39680 5360 39684
rect 5376 39740 5440 39744
rect 5376 39684 5380 39740
rect 5380 39684 5436 39740
rect 5436 39684 5440 39740
rect 5376 39680 5440 39684
rect 35856 39740 35920 39744
rect 35856 39684 35860 39740
rect 35860 39684 35916 39740
rect 35916 39684 35920 39740
rect 35856 39680 35920 39684
rect 35936 39740 36000 39744
rect 35936 39684 35940 39740
rect 35940 39684 35996 39740
rect 35996 39684 36000 39740
rect 35936 39680 36000 39684
rect 36016 39740 36080 39744
rect 36016 39684 36020 39740
rect 36020 39684 36076 39740
rect 36076 39684 36080 39740
rect 36016 39680 36080 39684
rect 36096 39740 36160 39744
rect 36096 39684 36100 39740
rect 36100 39684 36156 39740
rect 36156 39684 36160 39740
rect 36096 39680 36160 39684
rect 66576 39740 66640 39744
rect 66576 39684 66580 39740
rect 66580 39684 66636 39740
rect 66636 39684 66640 39740
rect 66576 39680 66640 39684
rect 66656 39740 66720 39744
rect 66656 39684 66660 39740
rect 66660 39684 66716 39740
rect 66716 39684 66720 39740
rect 66656 39680 66720 39684
rect 66736 39740 66800 39744
rect 66736 39684 66740 39740
rect 66740 39684 66796 39740
rect 66796 39684 66800 39740
rect 66736 39680 66800 39684
rect 66816 39740 66880 39744
rect 66816 39684 66820 39740
rect 66820 39684 66876 39740
rect 66876 39684 66880 39740
rect 66816 39680 66880 39684
rect 5796 39196 5860 39200
rect 5796 39140 5800 39196
rect 5800 39140 5856 39196
rect 5856 39140 5860 39196
rect 5796 39136 5860 39140
rect 5876 39196 5940 39200
rect 5876 39140 5880 39196
rect 5880 39140 5936 39196
rect 5936 39140 5940 39196
rect 5876 39136 5940 39140
rect 5956 39196 6020 39200
rect 5956 39140 5960 39196
rect 5960 39140 6016 39196
rect 6016 39140 6020 39196
rect 5956 39136 6020 39140
rect 6036 39196 6100 39200
rect 6036 39140 6040 39196
rect 6040 39140 6096 39196
rect 6096 39140 6100 39196
rect 6036 39136 6100 39140
rect 36516 39196 36580 39200
rect 36516 39140 36520 39196
rect 36520 39140 36576 39196
rect 36576 39140 36580 39196
rect 36516 39136 36580 39140
rect 36596 39196 36660 39200
rect 36596 39140 36600 39196
rect 36600 39140 36656 39196
rect 36656 39140 36660 39196
rect 36596 39136 36660 39140
rect 36676 39196 36740 39200
rect 36676 39140 36680 39196
rect 36680 39140 36736 39196
rect 36736 39140 36740 39196
rect 36676 39136 36740 39140
rect 36756 39196 36820 39200
rect 36756 39140 36760 39196
rect 36760 39140 36816 39196
rect 36816 39140 36820 39196
rect 36756 39136 36820 39140
rect 67236 39196 67300 39200
rect 67236 39140 67240 39196
rect 67240 39140 67296 39196
rect 67296 39140 67300 39196
rect 67236 39136 67300 39140
rect 67316 39196 67380 39200
rect 67316 39140 67320 39196
rect 67320 39140 67376 39196
rect 67376 39140 67380 39196
rect 67316 39136 67380 39140
rect 67396 39196 67460 39200
rect 67396 39140 67400 39196
rect 67400 39140 67456 39196
rect 67456 39140 67460 39196
rect 67396 39136 67460 39140
rect 67476 39196 67540 39200
rect 67476 39140 67480 39196
rect 67480 39140 67536 39196
rect 67536 39140 67540 39196
rect 67476 39136 67540 39140
rect 5136 38652 5200 38656
rect 5136 38596 5140 38652
rect 5140 38596 5196 38652
rect 5196 38596 5200 38652
rect 5136 38592 5200 38596
rect 5216 38652 5280 38656
rect 5216 38596 5220 38652
rect 5220 38596 5276 38652
rect 5276 38596 5280 38652
rect 5216 38592 5280 38596
rect 5296 38652 5360 38656
rect 5296 38596 5300 38652
rect 5300 38596 5356 38652
rect 5356 38596 5360 38652
rect 5296 38592 5360 38596
rect 5376 38652 5440 38656
rect 5376 38596 5380 38652
rect 5380 38596 5436 38652
rect 5436 38596 5440 38652
rect 5376 38592 5440 38596
rect 35856 38652 35920 38656
rect 35856 38596 35860 38652
rect 35860 38596 35916 38652
rect 35916 38596 35920 38652
rect 35856 38592 35920 38596
rect 35936 38652 36000 38656
rect 35936 38596 35940 38652
rect 35940 38596 35996 38652
rect 35996 38596 36000 38652
rect 35936 38592 36000 38596
rect 36016 38652 36080 38656
rect 36016 38596 36020 38652
rect 36020 38596 36076 38652
rect 36076 38596 36080 38652
rect 36016 38592 36080 38596
rect 36096 38652 36160 38656
rect 36096 38596 36100 38652
rect 36100 38596 36156 38652
rect 36156 38596 36160 38652
rect 36096 38592 36160 38596
rect 66576 38652 66640 38656
rect 66576 38596 66580 38652
rect 66580 38596 66636 38652
rect 66636 38596 66640 38652
rect 66576 38592 66640 38596
rect 66656 38652 66720 38656
rect 66656 38596 66660 38652
rect 66660 38596 66716 38652
rect 66716 38596 66720 38652
rect 66656 38592 66720 38596
rect 66736 38652 66800 38656
rect 66736 38596 66740 38652
rect 66740 38596 66796 38652
rect 66796 38596 66800 38652
rect 66736 38592 66800 38596
rect 66816 38652 66880 38656
rect 66816 38596 66820 38652
rect 66820 38596 66876 38652
rect 66876 38596 66880 38652
rect 66816 38592 66880 38596
rect 5796 38108 5860 38112
rect 5796 38052 5800 38108
rect 5800 38052 5856 38108
rect 5856 38052 5860 38108
rect 5796 38048 5860 38052
rect 5876 38108 5940 38112
rect 5876 38052 5880 38108
rect 5880 38052 5936 38108
rect 5936 38052 5940 38108
rect 5876 38048 5940 38052
rect 5956 38108 6020 38112
rect 5956 38052 5960 38108
rect 5960 38052 6016 38108
rect 6016 38052 6020 38108
rect 5956 38048 6020 38052
rect 6036 38108 6100 38112
rect 6036 38052 6040 38108
rect 6040 38052 6096 38108
rect 6096 38052 6100 38108
rect 6036 38048 6100 38052
rect 36516 38108 36580 38112
rect 36516 38052 36520 38108
rect 36520 38052 36576 38108
rect 36576 38052 36580 38108
rect 36516 38048 36580 38052
rect 36596 38108 36660 38112
rect 36596 38052 36600 38108
rect 36600 38052 36656 38108
rect 36656 38052 36660 38108
rect 36596 38048 36660 38052
rect 36676 38108 36740 38112
rect 36676 38052 36680 38108
rect 36680 38052 36736 38108
rect 36736 38052 36740 38108
rect 36676 38048 36740 38052
rect 36756 38108 36820 38112
rect 36756 38052 36760 38108
rect 36760 38052 36816 38108
rect 36816 38052 36820 38108
rect 36756 38048 36820 38052
rect 67236 38108 67300 38112
rect 67236 38052 67240 38108
rect 67240 38052 67296 38108
rect 67296 38052 67300 38108
rect 67236 38048 67300 38052
rect 67316 38108 67380 38112
rect 67316 38052 67320 38108
rect 67320 38052 67376 38108
rect 67376 38052 67380 38108
rect 67316 38048 67380 38052
rect 67396 38108 67460 38112
rect 67396 38052 67400 38108
rect 67400 38052 67456 38108
rect 67456 38052 67460 38108
rect 67396 38048 67460 38052
rect 67476 38108 67540 38112
rect 67476 38052 67480 38108
rect 67480 38052 67536 38108
rect 67536 38052 67540 38108
rect 67476 38048 67540 38052
rect 5136 37564 5200 37568
rect 5136 37508 5140 37564
rect 5140 37508 5196 37564
rect 5196 37508 5200 37564
rect 5136 37504 5200 37508
rect 5216 37564 5280 37568
rect 5216 37508 5220 37564
rect 5220 37508 5276 37564
rect 5276 37508 5280 37564
rect 5216 37504 5280 37508
rect 5296 37564 5360 37568
rect 5296 37508 5300 37564
rect 5300 37508 5356 37564
rect 5356 37508 5360 37564
rect 5296 37504 5360 37508
rect 5376 37564 5440 37568
rect 5376 37508 5380 37564
rect 5380 37508 5436 37564
rect 5436 37508 5440 37564
rect 5376 37504 5440 37508
rect 35856 37564 35920 37568
rect 35856 37508 35860 37564
rect 35860 37508 35916 37564
rect 35916 37508 35920 37564
rect 35856 37504 35920 37508
rect 35936 37564 36000 37568
rect 35936 37508 35940 37564
rect 35940 37508 35996 37564
rect 35996 37508 36000 37564
rect 35936 37504 36000 37508
rect 36016 37564 36080 37568
rect 36016 37508 36020 37564
rect 36020 37508 36076 37564
rect 36076 37508 36080 37564
rect 36016 37504 36080 37508
rect 36096 37564 36160 37568
rect 36096 37508 36100 37564
rect 36100 37508 36156 37564
rect 36156 37508 36160 37564
rect 36096 37504 36160 37508
rect 66576 37564 66640 37568
rect 66576 37508 66580 37564
rect 66580 37508 66636 37564
rect 66636 37508 66640 37564
rect 66576 37504 66640 37508
rect 66656 37564 66720 37568
rect 66656 37508 66660 37564
rect 66660 37508 66716 37564
rect 66716 37508 66720 37564
rect 66656 37504 66720 37508
rect 66736 37564 66800 37568
rect 66736 37508 66740 37564
rect 66740 37508 66796 37564
rect 66796 37508 66800 37564
rect 66736 37504 66800 37508
rect 66816 37564 66880 37568
rect 66816 37508 66820 37564
rect 66820 37508 66876 37564
rect 66876 37508 66880 37564
rect 66816 37504 66880 37508
rect 5796 37020 5860 37024
rect 5796 36964 5800 37020
rect 5800 36964 5856 37020
rect 5856 36964 5860 37020
rect 5796 36960 5860 36964
rect 5876 37020 5940 37024
rect 5876 36964 5880 37020
rect 5880 36964 5936 37020
rect 5936 36964 5940 37020
rect 5876 36960 5940 36964
rect 5956 37020 6020 37024
rect 5956 36964 5960 37020
rect 5960 36964 6016 37020
rect 6016 36964 6020 37020
rect 5956 36960 6020 36964
rect 6036 37020 6100 37024
rect 6036 36964 6040 37020
rect 6040 36964 6096 37020
rect 6096 36964 6100 37020
rect 6036 36960 6100 36964
rect 36516 37020 36580 37024
rect 36516 36964 36520 37020
rect 36520 36964 36576 37020
rect 36576 36964 36580 37020
rect 36516 36960 36580 36964
rect 36596 37020 36660 37024
rect 36596 36964 36600 37020
rect 36600 36964 36656 37020
rect 36656 36964 36660 37020
rect 36596 36960 36660 36964
rect 36676 37020 36740 37024
rect 36676 36964 36680 37020
rect 36680 36964 36736 37020
rect 36736 36964 36740 37020
rect 36676 36960 36740 36964
rect 36756 37020 36820 37024
rect 36756 36964 36760 37020
rect 36760 36964 36816 37020
rect 36816 36964 36820 37020
rect 36756 36960 36820 36964
rect 67236 37020 67300 37024
rect 67236 36964 67240 37020
rect 67240 36964 67296 37020
rect 67296 36964 67300 37020
rect 67236 36960 67300 36964
rect 67316 37020 67380 37024
rect 67316 36964 67320 37020
rect 67320 36964 67376 37020
rect 67376 36964 67380 37020
rect 67316 36960 67380 36964
rect 67396 37020 67460 37024
rect 67396 36964 67400 37020
rect 67400 36964 67456 37020
rect 67456 36964 67460 37020
rect 67396 36960 67460 36964
rect 67476 37020 67540 37024
rect 67476 36964 67480 37020
rect 67480 36964 67536 37020
rect 67536 36964 67540 37020
rect 67476 36960 67540 36964
rect 5136 36476 5200 36480
rect 5136 36420 5140 36476
rect 5140 36420 5196 36476
rect 5196 36420 5200 36476
rect 5136 36416 5200 36420
rect 5216 36476 5280 36480
rect 5216 36420 5220 36476
rect 5220 36420 5276 36476
rect 5276 36420 5280 36476
rect 5216 36416 5280 36420
rect 5296 36476 5360 36480
rect 5296 36420 5300 36476
rect 5300 36420 5356 36476
rect 5356 36420 5360 36476
rect 5296 36416 5360 36420
rect 5376 36476 5440 36480
rect 5376 36420 5380 36476
rect 5380 36420 5436 36476
rect 5436 36420 5440 36476
rect 5376 36416 5440 36420
rect 35856 36476 35920 36480
rect 35856 36420 35860 36476
rect 35860 36420 35916 36476
rect 35916 36420 35920 36476
rect 35856 36416 35920 36420
rect 35936 36476 36000 36480
rect 35936 36420 35940 36476
rect 35940 36420 35996 36476
rect 35996 36420 36000 36476
rect 35936 36416 36000 36420
rect 36016 36476 36080 36480
rect 36016 36420 36020 36476
rect 36020 36420 36076 36476
rect 36076 36420 36080 36476
rect 36016 36416 36080 36420
rect 36096 36476 36160 36480
rect 36096 36420 36100 36476
rect 36100 36420 36156 36476
rect 36156 36420 36160 36476
rect 36096 36416 36160 36420
rect 66576 36476 66640 36480
rect 66576 36420 66580 36476
rect 66580 36420 66636 36476
rect 66636 36420 66640 36476
rect 66576 36416 66640 36420
rect 66656 36476 66720 36480
rect 66656 36420 66660 36476
rect 66660 36420 66716 36476
rect 66716 36420 66720 36476
rect 66656 36416 66720 36420
rect 66736 36476 66800 36480
rect 66736 36420 66740 36476
rect 66740 36420 66796 36476
rect 66796 36420 66800 36476
rect 66736 36416 66800 36420
rect 66816 36476 66880 36480
rect 66816 36420 66820 36476
rect 66820 36420 66876 36476
rect 66876 36420 66880 36476
rect 66816 36416 66880 36420
rect 5796 35932 5860 35936
rect 5796 35876 5800 35932
rect 5800 35876 5856 35932
rect 5856 35876 5860 35932
rect 5796 35872 5860 35876
rect 5876 35932 5940 35936
rect 5876 35876 5880 35932
rect 5880 35876 5936 35932
rect 5936 35876 5940 35932
rect 5876 35872 5940 35876
rect 5956 35932 6020 35936
rect 5956 35876 5960 35932
rect 5960 35876 6016 35932
rect 6016 35876 6020 35932
rect 5956 35872 6020 35876
rect 6036 35932 6100 35936
rect 6036 35876 6040 35932
rect 6040 35876 6096 35932
rect 6096 35876 6100 35932
rect 6036 35872 6100 35876
rect 36516 35932 36580 35936
rect 36516 35876 36520 35932
rect 36520 35876 36576 35932
rect 36576 35876 36580 35932
rect 36516 35872 36580 35876
rect 36596 35932 36660 35936
rect 36596 35876 36600 35932
rect 36600 35876 36656 35932
rect 36656 35876 36660 35932
rect 36596 35872 36660 35876
rect 36676 35932 36740 35936
rect 36676 35876 36680 35932
rect 36680 35876 36736 35932
rect 36736 35876 36740 35932
rect 36676 35872 36740 35876
rect 36756 35932 36820 35936
rect 36756 35876 36760 35932
rect 36760 35876 36816 35932
rect 36816 35876 36820 35932
rect 36756 35872 36820 35876
rect 67236 35932 67300 35936
rect 67236 35876 67240 35932
rect 67240 35876 67296 35932
rect 67296 35876 67300 35932
rect 67236 35872 67300 35876
rect 67316 35932 67380 35936
rect 67316 35876 67320 35932
rect 67320 35876 67376 35932
rect 67376 35876 67380 35932
rect 67316 35872 67380 35876
rect 67396 35932 67460 35936
rect 67396 35876 67400 35932
rect 67400 35876 67456 35932
rect 67456 35876 67460 35932
rect 67396 35872 67460 35876
rect 67476 35932 67540 35936
rect 67476 35876 67480 35932
rect 67480 35876 67536 35932
rect 67536 35876 67540 35932
rect 67476 35872 67540 35876
rect 5136 35388 5200 35392
rect 5136 35332 5140 35388
rect 5140 35332 5196 35388
rect 5196 35332 5200 35388
rect 5136 35328 5200 35332
rect 5216 35388 5280 35392
rect 5216 35332 5220 35388
rect 5220 35332 5276 35388
rect 5276 35332 5280 35388
rect 5216 35328 5280 35332
rect 5296 35388 5360 35392
rect 5296 35332 5300 35388
rect 5300 35332 5356 35388
rect 5356 35332 5360 35388
rect 5296 35328 5360 35332
rect 5376 35388 5440 35392
rect 5376 35332 5380 35388
rect 5380 35332 5436 35388
rect 5436 35332 5440 35388
rect 5376 35328 5440 35332
rect 35856 35388 35920 35392
rect 35856 35332 35860 35388
rect 35860 35332 35916 35388
rect 35916 35332 35920 35388
rect 35856 35328 35920 35332
rect 35936 35388 36000 35392
rect 35936 35332 35940 35388
rect 35940 35332 35996 35388
rect 35996 35332 36000 35388
rect 35936 35328 36000 35332
rect 36016 35388 36080 35392
rect 36016 35332 36020 35388
rect 36020 35332 36076 35388
rect 36076 35332 36080 35388
rect 36016 35328 36080 35332
rect 36096 35388 36160 35392
rect 36096 35332 36100 35388
rect 36100 35332 36156 35388
rect 36156 35332 36160 35388
rect 36096 35328 36160 35332
rect 66576 35388 66640 35392
rect 66576 35332 66580 35388
rect 66580 35332 66636 35388
rect 66636 35332 66640 35388
rect 66576 35328 66640 35332
rect 66656 35388 66720 35392
rect 66656 35332 66660 35388
rect 66660 35332 66716 35388
rect 66716 35332 66720 35388
rect 66656 35328 66720 35332
rect 66736 35388 66800 35392
rect 66736 35332 66740 35388
rect 66740 35332 66796 35388
rect 66796 35332 66800 35388
rect 66736 35328 66800 35332
rect 66816 35388 66880 35392
rect 66816 35332 66820 35388
rect 66820 35332 66876 35388
rect 66876 35332 66880 35388
rect 66816 35328 66880 35332
rect 5796 34844 5860 34848
rect 5796 34788 5800 34844
rect 5800 34788 5856 34844
rect 5856 34788 5860 34844
rect 5796 34784 5860 34788
rect 5876 34844 5940 34848
rect 5876 34788 5880 34844
rect 5880 34788 5936 34844
rect 5936 34788 5940 34844
rect 5876 34784 5940 34788
rect 5956 34844 6020 34848
rect 5956 34788 5960 34844
rect 5960 34788 6016 34844
rect 6016 34788 6020 34844
rect 5956 34784 6020 34788
rect 6036 34844 6100 34848
rect 6036 34788 6040 34844
rect 6040 34788 6096 34844
rect 6096 34788 6100 34844
rect 6036 34784 6100 34788
rect 36516 34844 36580 34848
rect 36516 34788 36520 34844
rect 36520 34788 36576 34844
rect 36576 34788 36580 34844
rect 36516 34784 36580 34788
rect 36596 34844 36660 34848
rect 36596 34788 36600 34844
rect 36600 34788 36656 34844
rect 36656 34788 36660 34844
rect 36596 34784 36660 34788
rect 36676 34844 36740 34848
rect 36676 34788 36680 34844
rect 36680 34788 36736 34844
rect 36736 34788 36740 34844
rect 36676 34784 36740 34788
rect 36756 34844 36820 34848
rect 36756 34788 36760 34844
rect 36760 34788 36816 34844
rect 36816 34788 36820 34844
rect 36756 34784 36820 34788
rect 67236 34844 67300 34848
rect 67236 34788 67240 34844
rect 67240 34788 67296 34844
rect 67296 34788 67300 34844
rect 67236 34784 67300 34788
rect 67316 34844 67380 34848
rect 67316 34788 67320 34844
rect 67320 34788 67376 34844
rect 67376 34788 67380 34844
rect 67316 34784 67380 34788
rect 67396 34844 67460 34848
rect 67396 34788 67400 34844
rect 67400 34788 67456 34844
rect 67456 34788 67460 34844
rect 67396 34784 67460 34788
rect 67476 34844 67540 34848
rect 67476 34788 67480 34844
rect 67480 34788 67536 34844
rect 67536 34788 67540 34844
rect 67476 34784 67540 34788
rect 5136 34300 5200 34304
rect 5136 34244 5140 34300
rect 5140 34244 5196 34300
rect 5196 34244 5200 34300
rect 5136 34240 5200 34244
rect 5216 34300 5280 34304
rect 5216 34244 5220 34300
rect 5220 34244 5276 34300
rect 5276 34244 5280 34300
rect 5216 34240 5280 34244
rect 5296 34300 5360 34304
rect 5296 34244 5300 34300
rect 5300 34244 5356 34300
rect 5356 34244 5360 34300
rect 5296 34240 5360 34244
rect 5376 34300 5440 34304
rect 5376 34244 5380 34300
rect 5380 34244 5436 34300
rect 5436 34244 5440 34300
rect 5376 34240 5440 34244
rect 35856 34300 35920 34304
rect 35856 34244 35860 34300
rect 35860 34244 35916 34300
rect 35916 34244 35920 34300
rect 35856 34240 35920 34244
rect 35936 34300 36000 34304
rect 35936 34244 35940 34300
rect 35940 34244 35996 34300
rect 35996 34244 36000 34300
rect 35936 34240 36000 34244
rect 36016 34300 36080 34304
rect 36016 34244 36020 34300
rect 36020 34244 36076 34300
rect 36076 34244 36080 34300
rect 36016 34240 36080 34244
rect 36096 34300 36160 34304
rect 36096 34244 36100 34300
rect 36100 34244 36156 34300
rect 36156 34244 36160 34300
rect 36096 34240 36160 34244
rect 66576 34300 66640 34304
rect 66576 34244 66580 34300
rect 66580 34244 66636 34300
rect 66636 34244 66640 34300
rect 66576 34240 66640 34244
rect 66656 34300 66720 34304
rect 66656 34244 66660 34300
rect 66660 34244 66716 34300
rect 66716 34244 66720 34300
rect 66656 34240 66720 34244
rect 66736 34300 66800 34304
rect 66736 34244 66740 34300
rect 66740 34244 66796 34300
rect 66796 34244 66800 34300
rect 66736 34240 66800 34244
rect 66816 34300 66880 34304
rect 66816 34244 66820 34300
rect 66820 34244 66876 34300
rect 66876 34244 66880 34300
rect 66816 34240 66880 34244
rect 5796 33756 5860 33760
rect 5796 33700 5800 33756
rect 5800 33700 5856 33756
rect 5856 33700 5860 33756
rect 5796 33696 5860 33700
rect 5876 33756 5940 33760
rect 5876 33700 5880 33756
rect 5880 33700 5936 33756
rect 5936 33700 5940 33756
rect 5876 33696 5940 33700
rect 5956 33756 6020 33760
rect 5956 33700 5960 33756
rect 5960 33700 6016 33756
rect 6016 33700 6020 33756
rect 5956 33696 6020 33700
rect 6036 33756 6100 33760
rect 6036 33700 6040 33756
rect 6040 33700 6096 33756
rect 6096 33700 6100 33756
rect 6036 33696 6100 33700
rect 36516 33756 36580 33760
rect 36516 33700 36520 33756
rect 36520 33700 36576 33756
rect 36576 33700 36580 33756
rect 36516 33696 36580 33700
rect 36596 33756 36660 33760
rect 36596 33700 36600 33756
rect 36600 33700 36656 33756
rect 36656 33700 36660 33756
rect 36596 33696 36660 33700
rect 36676 33756 36740 33760
rect 36676 33700 36680 33756
rect 36680 33700 36736 33756
rect 36736 33700 36740 33756
rect 36676 33696 36740 33700
rect 36756 33756 36820 33760
rect 36756 33700 36760 33756
rect 36760 33700 36816 33756
rect 36816 33700 36820 33756
rect 36756 33696 36820 33700
rect 67236 33756 67300 33760
rect 67236 33700 67240 33756
rect 67240 33700 67296 33756
rect 67296 33700 67300 33756
rect 67236 33696 67300 33700
rect 67316 33756 67380 33760
rect 67316 33700 67320 33756
rect 67320 33700 67376 33756
rect 67376 33700 67380 33756
rect 67316 33696 67380 33700
rect 67396 33756 67460 33760
rect 67396 33700 67400 33756
rect 67400 33700 67456 33756
rect 67456 33700 67460 33756
rect 67396 33696 67460 33700
rect 67476 33756 67540 33760
rect 67476 33700 67480 33756
rect 67480 33700 67536 33756
rect 67536 33700 67540 33756
rect 67476 33696 67540 33700
rect 5136 33212 5200 33216
rect 5136 33156 5140 33212
rect 5140 33156 5196 33212
rect 5196 33156 5200 33212
rect 5136 33152 5200 33156
rect 5216 33212 5280 33216
rect 5216 33156 5220 33212
rect 5220 33156 5276 33212
rect 5276 33156 5280 33212
rect 5216 33152 5280 33156
rect 5296 33212 5360 33216
rect 5296 33156 5300 33212
rect 5300 33156 5356 33212
rect 5356 33156 5360 33212
rect 5296 33152 5360 33156
rect 5376 33212 5440 33216
rect 5376 33156 5380 33212
rect 5380 33156 5436 33212
rect 5436 33156 5440 33212
rect 5376 33152 5440 33156
rect 35856 33212 35920 33216
rect 35856 33156 35860 33212
rect 35860 33156 35916 33212
rect 35916 33156 35920 33212
rect 35856 33152 35920 33156
rect 35936 33212 36000 33216
rect 35936 33156 35940 33212
rect 35940 33156 35996 33212
rect 35996 33156 36000 33212
rect 35936 33152 36000 33156
rect 36016 33212 36080 33216
rect 36016 33156 36020 33212
rect 36020 33156 36076 33212
rect 36076 33156 36080 33212
rect 36016 33152 36080 33156
rect 36096 33212 36160 33216
rect 36096 33156 36100 33212
rect 36100 33156 36156 33212
rect 36156 33156 36160 33212
rect 36096 33152 36160 33156
rect 66576 33212 66640 33216
rect 66576 33156 66580 33212
rect 66580 33156 66636 33212
rect 66636 33156 66640 33212
rect 66576 33152 66640 33156
rect 66656 33212 66720 33216
rect 66656 33156 66660 33212
rect 66660 33156 66716 33212
rect 66716 33156 66720 33212
rect 66656 33152 66720 33156
rect 66736 33212 66800 33216
rect 66736 33156 66740 33212
rect 66740 33156 66796 33212
rect 66796 33156 66800 33212
rect 66736 33152 66800 33156
rect 66816 33212 66880 33216
rect 66816 33156 66820 33212
rect 66820 33156 66876 33212
rect 66876 33156 66880 33212
rect 66816 33152 66880 33156
rect 5796 32668 5860 32672
rect 5796 32612 5800 32668
rect 5800 32612 5856 32668
rect 5856 32612 5860 32668
rect 5796 32608 5860 32612
rect 5876 32668 5940 32672
rect 5876 32612 5880 32668
rect 5880 32612 5936 32668
rect 5936 32612 5940 32668
rect 5876 32608 5940 32612
rect 5956 32668 6020 32672
rect 5956 32612 5960 32668
rect 5960 32612 6016 32668
rect 6016 32612 6020 32668
rect 5956 32608 6020 32612
rect 6036 32668 6100 32672
rect 6036 32612 6040 32668
rect 6040 32612 6096 32668
rect 6096 32612 6100 32668
rect 6036 32608 6100 32612
rect 36516 32668 36580 32672
rect 36516 32612 36520 32668
rect 36520 32612 36576 32668
rect 36576 32612 36580 32668
rect 36516 32608 36580 32612
rect 36596 32668 36660 32672
rect 36596 32612 36600 32668
rect 36600 32612 36656 32668
rect 36656 32612 36660 32668
rect 36596 32608 36660 32612
rect 36676 32668 36740 32672
rect 36676 32612 36680 32668
rect 36680 32612 36736 32668
rect 36736 32612 36740 32668
rect 36676 32608 36740 32612
rect 36756 32668 36820 32672
rect 36756 32612 36760 32668
rect 36760 32612 36816 32668
rect 36816 32612 36820 32668
rect 36756 32608 36820 32612
rect 67236 32668 67300 32672
rect 67236 32612 67240 32668
rect 67240 32612 67296 32668
rect 67296 32612 67300 32668
rect 67236 32608 67300 32612
rect 67316 32668 67380 32672
rect 67316 32612 67320 32668
rect 67320 32612 67376 32668
rect 67376 32612 67380 32668
rect 67316 32608 67380 32612
rect 67396 32668 67460 32672
rect 67396 32612 67400 32668
rect 67400 32612 67456 32668
rect 67456 32612 67460 32668
rect 67396 32608 67460 32612
rect 67476 32668 67540 32672
rect 67476 32612 67480 32668
rect 67480 32612 67536 32668
rect 67536 32612 67540 32668
rect 67476 32608 67540 32612
rect 5136 32124 5200 32128
rect 5136 32068 5140 32124
rect 5140 32068 5196 32124
rect 5196 32068 5200 32124
rect 5136 32064 5200 32068
rect 5216 32124 5280 32128
rect 5216 32068 5220 32124
rect 5220 32068 5276 32124
rect 5276 32068 5280 32124
rect 5216 32064 5280 32068
rect 5296 32124 5360 32128
rect 5296 32068 5300 32124
rect 5300 32068 5356 32124
rect 5356 32068 5360 32124
rect 5296 32064 5360 32068
rect 5376 32124 5440 32128
rect 5376 32068 5380 32124
rect 5380 32068 5436 32124
rect 5436 32068 5440 32124
rect 5376 32064 5440 32068
rect 35856 32124 35920 32128
rect 35856 32068 35860 32124
rect 35860 32068 35916 32124
rect 35916 32068 35920 32124
rect 35856 32064 35920 32068
rect 35936 32124 36000 32128
rect 35936 32068 35940 32124
rect 35940 32068 35996 32124
rect 35996 32068 36000 32124
rect 35936 32064 36000 32068
rect 36016 32124 36080 32128
rect 36016 32068 36020 32124
rect 36020 32068 36076 32124
rect 36076 32068 36080 32124
rect 36016 32064 36080 32068
rect 36096 32124 36160 32128
rect 36096 32068 36100 32124
rect 36100 32068 36156 32124
rect 36156 32068 36160 32124
rect 36096 32064 36160 32068
rect 66576 32124 66640 32128
rect 66576 32068 66580 32124
rect 66580 32068 66636 32124
rect 66636 32068 66640 32124
rect 66576 32064 66640 32068
rect 66656 32124 66720 32128
rect 66656 32068 66660 32124
rect 66660 32068 66716 32124
rect 66716 32068 66720 32124
rect 66656 32064 66720 32068
rect 66736 32124 66800 32128
rect 66736 32068 66740 32124
rect 66740 32068 66796 32124
rect 66796 32068 66800 32124
rect 66736 32064 66800 32068
rect 66816 32124 66880 32128
rect 66816 32068 66820 32124
rect 66820 32068 66876 32124
rect 66876 32068 66880 32124
rect 66816 32064 66880 32068
rect 5796 31580 5860 31584
rect 5796 31524 5800 31580
rect 5800 31524 5856 31580
rect 5856 31524 5860 31580
rect 5796 31520 5860 31524
rect 5876 31580 5940 31584
rect 5876 31524 5880 31580
rect 5880 31524 5936 31580
rect 5936 31524 5940 31580
rect 5876 31520 5940 31524
rect 5956 31580 6020 31584
rect 5956 31524 5960 31580
rect 5960 31524 6016 31580
rect 6016 31524 6020 31580
rect 5956 31520 6020 31524
rect 6036 31580 6100 31584
rect 6036 31524 6040 31580
rect 6040 31524 6096 31580
rect 6096 31524 6100 31580
rect 6036 31520 6100 31524
rect 36516 31580 36580 31584
rect 36516 31524 36520 31580
rect 36520 31524 36576 31580
rect 36576 31524 36580 31580
rect 36516 31520 36580 31524
rect 36596 31580 36660 31584
rect 36596 31524 36600 31580
rect 36600 31524 36656 31580
rect 36656 31524 36660 31580
rect 36596 31520 36660 31524
rect 36676 31580 36740 31584
rect 36676 31524 36680 31580
rect 36680 31524 36736 31580
rect 36736 31524 36740 31580
rect 36676 31520 36740 31524
rect 36756 31580 36820 31584
rect 36756 31524 36760 31580
rect 36760 31524 36816 31580
rect 36816 31524 36820 31580
rect 36756 31520 36820 31524
rect 67236 31580 67300 31584
rect 67236 31524 67240 31580
rect 67240 31524 67296 31580
rect 67296 31524 67300 31580
rect 67236 31520 67300 31524
rect 67316 31580 67380 31584
rect 67316 31524 67320 31580
rect 67320 31524 67376 31580
rect 67376 31524 67380 31580
rect 67316 31520 67380 31524
rect 67396 31580 67460 31584
rect 67396 31524 67400 31580
rect 67400 31524 67456 31580
rect 67456 31524 67460 31580
rect 67396 31520 67460 31524
rect 67476 31580 67540 31584
rect 67476 31524 67480 31580
rect 67480 31524 67536 31580
rect 67536 31524 67540 31580
rect 67476 31520 67540 31524
rect 5136 31036 5200 31040
rect 5136 30980 5140 31036
rect 5140 30980 5196 31036
rect 5196 30980 5200 31036
rect 5136 30976 5200 30980
rect 5216 31036 5280 31040
rect 5216 30980 5220 31036
rect 5220 30980 5276 31036
rect 5276 30980 5280 31036
rect 5216 30976 5280 30980
rect 5296 31036 5360 31040
rect 5296 30980 5300 31036
rect 5300 30980 5356 31036
rect 5356 30980 5360 31036
rect 5296 30976 5360 30980
rect 5376 31036 5440 31040
rect 5376 30980 5380 31036
rect 5380 30980 5436 31036
rect 5436 30980 5440 31036
rect 5376 30976 5440 30980
rect 35856 31036 35920 31040
rect 35856 30980 35860 31036
rect 35860 30980 35916 31036
rect 35916 30980 35920 31036
rect 35856 30976 35920 30980
rect 35936 31036 36000 31040
rect 35936 30980 35940 31036
rect 35940 30980 35996 31036
rect 35996 30980 36000 31036
rect 35936 30976 36000 30980
rect 36016 31036 36080 31040
rect 36016 30980 36020 31036
rect 36020 30980 36076 31036
rect 36076 30980 36080 31036
rect 36016 30976 36080 30980
rect 36096 31036 36160 31040
rect 36096 30980 36100 31036
rect 36100 30980 36156 31036
rect 36156 30980 36160 31036
rect 36096 30976 36160 30980
rect 66576 31036 66640 31040
rect 66576 30980 66580 31036
rect 66580 30980 66636 31036
rect 66636 30980 66640 31036
rect 66576 30976 66640 30980
rect 66656 31036 66720 31040
rect 66656 30980 66660 31036
rect 66660 30980 66716 31036
rect 66716 30980 66720 31036
rect 66656 30976 66720 30980
rect 66736 31036 66800 31040
rect 66736 30980 66740 31036
rect 66740 30980 66796 31036
rect 66796 30980 66800 31036
rect 66736 30976 66800 30980
rect 66816 31036 66880 31040
rect 66816 30980 66820 31036
rect 66820 30980 66876 31036
rect 66876 30980 66880 31036
rect 66816 30976 66880 30980
rect 5796 30492 5860 30496
rect 5796 30436 5800 30492
rect 5800 30436 5856 30492
rect 5856 30436 5860 30492
rect 5796 30432 5860 30436
rect 5876 30492 5940 30496
rect 5876 30436 5880 30492
rect 5880 30436 5936 30492
rect 5936 30436 5940 30492
rect 5876 30432 5940 30436
rect 5956 30492 6020 30496
rect 5956 30436 5960 30492
rect 5960 30436 6016 30492
rect 6016 30436 6020 30492
rect 5956 30432 6020 30436
rect 6036 30492 6100 30496
rect 6036 30436 6040 30492
rect 6040 30436 6096 30492
rect 6096 30436 6100 30492
rect 6036 30432 6100 30436
rect 36516 30492 36580 30496
rect 36516 30436 36520 30492
rect 36520 30436 36576 30492
rect 36576 30436 36580 30492
rect 36516 30432 36580 30436
rect 36596 30492 36660 30496
rect 36596 30436 36600 30492
rect 36600 30436 36656 30492
rect 36656 30436 36660 30492
rect 36596 30432 36660 30436
rect 36676 30492 36740 30496
rect 36676 30436 36680 30492
rect 36680 30436 36736 30492
rect 36736 30436 36740 30492
rect 36676 30432 36740 30436
rect 36756 30492 36820 30496
rect 36756 30436 36760 30492
rect 36760 30436 36816 30492
rect 36816 30436 36820 30492
rect 36756 30432 36820 30436
rect 67236 30492 67300 30496
rect 67236 30436 67240 30492
rect 67240 30436 67296 30492
rect 67296 30436 67300 30492
rect 67236 30432 67300 30436
rect 67316 30492 67380 30496
rect 67316 30436 67320 30492
rect 67320 30436 67376 30492
rect 67376 30436 67380 30492
rect 67316 30432 67380 30436
rect 67396 30492 67460 30496
rect 67396 30436 67400 30492
rect 67400 30436 67456 30492
rect 67456 30436 67460 30492
rect 67396 30432 67460 30436
rect 67476 30492 67540 30496
rect 67476 30436 67480 30492
rect 67480 30436 67536 30492
rect 67536 30436 67540 30492
rect 67476 30432 67540 30436
rect 5136 29948 5200 29952
rect 5136 29892 5140 29948
rect 5140 29892 5196 29948
rect 5196 29892 5200 29948
rect 5136 29888 5200 29892
rect 5216 29948 5280 29952
rect 5216 29892 5220 29948
rect 5220 29892 5276 29948
rect 5276 29892 5280 29948
rect 5216 29888 5280 29892
rect 5296 29948 5360 29952
rect 5296 29892 5300 29948
rect 5300 29892 5356 29948
rect 5356 29892 5360 29948
rect 5296 29888 5360 29892
rect 5376 29948 5440 29952
rect 5376 29892 5380 29948
rect 5380 29892 5436 29948
rect 5436 29892 5440 29948
rect 5376 29888 5440 29892
rect 35856 29948 35920 29952
rect 35856 29892 35860 29948
rect 35860 29892 35916 29948
rect 35916 29892 35920 29948
rect 35856 29888 35920 29892
rect 35936 29948 36000 29952
rect 35936 29892 35940 29948
rect 35940 29892 35996 29948
rect 35996 29892 36000 29948
rect 35936 29888 36000 29892
rect 36016 29948 36080 29952
rect 36016 29892 36020 29948
rect 36020 29892 36076 29948
rect 36076 29892 36080 29948
rect 36016 29888 36080 29892
rect 36096 29948 36160 29952
rect 36096 29892 36100 29948
rect 36100 29892 36156 29948
rect 36156 29892 36160 29948
rect 36096 29888 36160 29892
rect 66576 29948 66640 29952
rect 66576 29892 66580 29948
rect 66580 29892 66636 29948
rect 66636 29892 66640 29948
rect 66576 29888 66640 29892
rect 66656 29948 66720 29952
rect 66656 29892 66660 29948
rect 66660 29892 66716 29948
rect 66716 29892 66720 29948
rect 66656 29888 66720 29892
rect 66736 29948 66800 29952
rect 66736 29892 66740 29948
rect 66740 29892 66796 29948
rect 66796 29892 66800 29948
rect 66736 29888 66800 29892
rect 66816 29948 66880 29952
rect 66816 29892 66820 29948
rect 66820 29892 66876 29948
rect 66876 29892 66880 29948
rect 66816 29888 66880 29892
rect 5796 29404 5860 29408
rect 5796 29348 5800 29404
rect 5800 29348 5856 29404
rect 5856 29348 5860 29404
rect 5796 29344 5860 29348
rect 5876 29404 5940 29408
rect 5876 29348 5880 29404
rect 5880 29348 5936 29404
rect 5936 29348 5940 29404
rect 5876 29344 5940 29348
rect 5956 29404 6020 29408
rect 5956 29348 5960 29404
rect 5960 29348 6016 29404
rect 6016 29348 6020 29404
rect 5956 29344 6020 29348
rect 6036 29404 6100 29408
rect 6036 29348 6040 29404
rect 6040 29348 6096 29404
rect 6096 29348 6100 29404
rect 6036 29344 6100 29348
rect 36516 29404 36580 29408
rect 36516 29348 36520 29404
rect 36520 29348 36576 29404
rect 36576 29348 36580 29404
rect 36516 29344 36580 29348
rect 36596 29404 36660 29408
rect 36596 29348 36600 29404
rect 36600 29348 36656 29404
rect 36656 29348 36660 29404
rect 36596 29344 36660 29348
rect 36676 29404 36740 29408
rect 36676 29348 36680 29404
rect 36680 29348 36736 29404
rect 36736 29348 36740 29404
rect 36676 29344 36740 29348
rect 36756 29404 36820 29408
rect 36756 29348 36760 29404
rect 36760 29348 36816 29404
rect 36816 29348 36820 29404
rect 36756 29344 36820 29348
rect 67236 29404 67300 29408
rect 67236 29348 67240 29404
rect 67240 29348 67296 29404
rect 67296 29348 67300 29404
rect 67236 29344 67300 29348
rect 67316 29404 67380 29408
rect 67316 29348 67320 29404
rect 67320 29348 67376 29404
rect 67376 29348 67380 29404
rect 67316 29344 67380 29348
rect 67396 29404 67460 29408
rect 67396 29348 67400 29404
rect 67400 29348 67456 29404
rect 67456 29348 67460 29404
rect 67396 29344 67460 29348
rect 67476 29404 67540 29408
rect 67476 29348 67480 29404
rect 67480 29348 67536 29404
rect 67536 29348 67540 29404
rect 67476 29344 67540 29348
rect 5136 28860 5200 28864
rect 5136 28804 5140 28860
rect 5140 28804 5196 28860
rect 5196 28804 5200 28860
rect 5136 28800 5200 28804
rect 5216 28860 5280 28864
rect 5216 28804 5220 28860
rect 5220 28804 5276 28860
rect 5276 28804 5280 28860
rect 5216 28800 5280 28804
rect 5296 28860 5360 28864
rect 5296 28804 5300 28860
rect 5300 28804 5356 28860
rect 5356 28804 5360 28860
rect 5296 28800 5360 28804
rect 5376 28860 5440 28864
rect 5376 28804 5380 28860
rect 5380 28804 5436 28860
rect 5436 28804 5440 28860
rect 5376 28800 5440 28804
rect 35856 28860 35920 28864
rect 35856 28804 35860 28860
rect 35860 28804 35916 28860
rect 35916 28804 35920 28860
rect 35856 28800 35920 28804
rect 35936 28860 36000 28864
rect 35936 28804 35940 28860
rect 35940 28804 35996 28860
rect 35996 28804 36000 28860
rect 35936 28800 36000 28804
rect 36016 28860 36080 28864
rect 36016 28804 36020 28860
rect 36020 28804 36076 28860
rect 36076 28804 36080 28860
rect 36016 28800 36080 28804
rect 36096 28860 36160 28864
rect 36096 28804 36100 28860
rect 36100 28804 36156 28860
rect 36156 28804 36160 28860
rect 36096 28800 36160 28804
rect 66576 28860 66640 28864
rect 66576 28804 66580 28860
rect 66580 28804 66636 28860
rect 66636 28804 66640 28860
rect 66576 28800 66640 28804
rect 66656 28860 66720 28864
rect 66656 28804 66660 28860
rect 66660 28804 66716 28860
rect 66716 28804 66720 28860
rect 66656 28800 66720 28804
rect 66736 28860 66800 28864
rect 66736 28804 66740 28860
rect 66740 28804 66796 28860
rect 66796 28804 66800 28860
rect 66736 28800 66800 28804
rect 66816 28860 66880 28864
rect 66816 28804 66820 28860
rect 66820 28804 66876 28860
rect 66876 28804 66880 28860
rect 66816 28800 66880 28804
rect 5796 28316 5860 28320
rect 5796 28260 5800 28316
rect 5800 28260 5856 28316
rect 5856 28260 5860 28316
rect 5796 28256 5860 28260
rect 5876 28316 5940 28320
rect 5876 28260 5880 28316
rect 5880 28260 5936 28316
rect 5936 28260 5940 28316
rect 5876 28256 5940 28260
rect 5956 28316 6020 28320
rect 5956 28260 5960 28316
rect 5960 28260 6016 28316
rect 6016 28260 6020 28316
rect 5956 28256 6020 28260
rect 6036 28316 6100 28320
rect 6036 28260 6040 28316
rect 6040 28260 6096 28316
rect 6096 28260 6100 28316
rect 6036 28256 6100 28260
rect 36516 28316 36580 28320
rect 36516 28260 36520 28316
rect 36520 28260 36576 28316
rect 36576 28260 36580 28316
rect 36516 28256 36580 28260
rect 36596 28316 36660 28320
rect 36596 28260 36600 28316
rect 36600 28260 36656 28316
rect 36656 28260 36660 28316
rect 36596 28256 36660 28260
rect 36676 28316 36740 28320
rect 36676 28260 36680 28316
rect 36680 28260 36736 28316
rect 36736 28260 36740 28316
rect 36676 28256 36740 28260
rect 36756 28316 36820 28320
rect 36756 28260 36760 28316
rect 36760 28260 36816 28316
rect 36816 28260 36820 28316
rect 36756 28256 36820 28260
rect 67236 28316 67300 28320
rect 67236 28260 67240 28316
rect 67240 28260 67296 28316
rect 67296 28260 67300 28316
rect 67236 28256 67300 28260
rect 67316 28316 67380 28320
rect 67316 28260 67320 28316
rect 67320 28260 67376 28316
rect 67376 28260 67380 28316
rect 67316 28256 67380 28260
rect 67396 28316 67460 28320
rect 67396 28260 67400 28316
rect 67400 28260 67456 28316
rect 67456 28260 67460 28316
rect 67396 28256 67460 28260
rect 67476 28316 67540 28320
rect 67476 28260 67480 28316
rect 67480 28260 67536 28316
rect 67536 28260 67540 28316
rect 67476 28256 67540 28260
rect 5136 27772 5200 27776
rect 5136 27716 5140 27772
rect 5140 27716 5196 27772
rect 5196 27716 5200 27772
rect 5136 27712 5200 27716
rect 5216 27772 5280 27776
rect 5216 27716 5220 27772
rect 5220 27716 5276 27772
rect 5276 27716 5280 27772
rect 5216 27712 5280 27716
rect 5296 27772 5360 27776
rect 5296 27716 5300 27772
rect 5300 27716 5356 27772
rect 5356 27716 5360 27772
rect 5296 27712 5360 27716
rect 5376 27772 5440 27776
rect 5376 27716 5380 27772
rect 5380 27716 5436 27772
rect 5436 27716 5440 27772
rect 5376 27712 5440 27716
rect 35856 27772 35920 27776
rect 35856 27716 35860 27772
rect 35860 27716 35916 27772
rect 35916 27716 35920 27772
rect 35856 27712 35920 27716
rect 35936 27772 36000 27776
rect 35936 27716 35940 27772
rect 35940 27716 35996 27772
rect 35996 27716 36000 27772
rect 35936 27712 36000 27716
rect 36016 27772 36080 27776
rect 36016 27716 36020 27772
rect 36020 27716 36076 27772
rect 36076 27716 36080 27772
rect 36016 27712 36080 27716
rect 36096 27772 36160 27776
rect 36096 27716 36100 27772
rect 36100 27716 36156 27772
rect 36156 27716 36160 27772
rect 36096 27712 36160 27716
rect 66576 27772 66640 27776
rect 66576 27716 66580 27772
rect 66580 27716 66636 27772
rect 66636 27716 66640 27772
rect 66576 27712 66640 27716
rect 66656 27772 66720 27776
rect 66656 27716 66660 27772
rect 66660 27716 66716 27772
rect 66716 27716 66720 27772
rect 66656 27712 66720 27716
rect 66736 27772 66800 27776
rect 66736 27716 66740 27772
rect 66740 27716 66796 27772
rect 66796 27716 66800 27772
rect 66736 27712 66800 27716
rect 66816 27772 66880 27776
rect 66816 27716 66820 27772
rect 66820 27716 66876 27772
rect 66876 27716 66880 27772
rect 66816 27712 66880 27716
rect 5796 27228 5860 27232
rect 5796 27172 5800 27228
rect 5800 27172 5856 27228
rect 5856 27172 5860 27228
rect 5796 27168 5860 27172
rect 5876 27228 5940 27232
rect 5876 27172 5880 27228
rect 5880 27172 5936 27228
rect 5936 27172 5940 27228
rect 5876 27168 5940 27172
rect 5956 27228 6020 27232
rect 5956 27172 5960 27228
rect 5960 27172 6016 27228
rect 6016 27172 6020 27228
rect 5956 27168 6020 27172
rect 6036 27228 6100 27232
rect 6036 27172 6040 27228
rect 6040 27172 6096 27228
rect 6096 27172 6100 27228
rect 6036 27168 6100 27172
rect 36516 27228 36580 27232
rect 36516 27172 36520 27228
rect 36520 27172 36576 27228
rect 36576 27172 36580 27228
rect 36516 27168 36580 27172
rect 36596 27228 36660 27232
rect 36596 27172 36600 27228
rect 36600 27172 36656 27228
rect 36656 27172 36660 27228
rect 36596 27168 36660 27172
rect 36676 27228 36740 27232
rect 36676 27172 36680 27228
rect 36680 27172 36736 27228
rect 36736 27172 36740 27228
rect 36676 27168 36740 27172
rect 36756 27228 36820 27232
rect 36756 27172 36760 27228
rect 36760 27172 36816 27228
rect 36816 27172 36820 27228
rect 36756 27168 36820 27172
rect 67236 27228 67300 27232
rect 67236 27172 67240 27228
rect 67240 27172 67296 27228
rect 67296 27172 67300 27228
rect 67236 27168 67300 27172
rect 67316 27228 67380 27232
rect 67316 27172 67320 27228
rect 67320 27172 67376 27228
rect 67376 27172 67380 27228
rect 67316 27168 67380 27172
rect 67396 27228 67460 27232
rect 67396 27172 67400 27228
rect 67400 27172 67456 27228
rect 67456 27172 67460 27228
rect 67396 27168 67460 27172
rect 67476 27228 67540 27232
rect 67476 27172 67480 27228
rect 67480 27172 67536 27228
rect 67536 27172 67540 27228
rect 67476 27168 67540 27172
rect 5136 26684 5200 26688
rect 5136 26628 5140 26684
rect 5140 26628 5196 26684
rect 5196 26628 5200 26684
rect 5136 26624 5200 26628
rect 5216 26684 5280 26688
rect 5216 26628 5220 26684
rect 5220 26628 5276 26684
rect 5276 26628 5280 26684
rect 5216 26624 5280 26628
rect 5296 26684 5360 26688
rect 5296 26628 5300 26684
rect 5300 26628 5356 26684
rect 5356 26628 5360 26684
rect 5296 26624 5360 26628
rect 5376 26684 5440 26688
rect 5376 26628 5380 26684
rect 5380 26628 5436 26684
rect 5436 26628 5440 26684
rect 5376 26624 5440 26628
rect 35856 26684 35920 26688
rect 35856 26628 35860 26684
rect 35860 26628 35916 26684
rect 35916 26628 35920 26684
rect 35856 26624 35920 26628
rect 35936 26684 36000 26688
rect 35936 26628 35940 26684
rect 35940 26628 35996 26684
rect 35996 26628 36000 26684
rect 35936 26624 36000 26628
rect 36016 26684 36080 26688
rect 36016 26628 36020 26684
rect 36020 26628 36076 26684
rect 36076 26628 36080 26684
rect 36016 26624 36080 26628
rect 36096 26684 36160 26688
rect 36096 26628 36100 26684
rect 36100 26628 36156 26684
rect 36156 26628 36160 26684
rect 36096 26624 36160 26628
rect 66576 26684 66640 26688
rect 66576 26628 66580 26684
rect 66580 26628 66636 26684
rect 66636 26628 66640 26684
rect 66576 26624 66640 26628
rect 66656 26684 66720 26688
rect 66656 26628 66660 26684
rect 66660 26628 66716 26684
rect 66716 26628 66720 26684
rect 66656 26624 66720 26628
rect 66736 26684 66800 26688
rect 66736 26628 66740 26684
rect 66740 26628 66796 26684
rect 66796 26628 66800 26684
rect 66736 26624 66800 26628
rect 66816 26684 66880 26688
rect 66816 26628 66820 26684
rect 66820 26628 66876 26684
rect 66876 26628 66880 26684
rect 66816 26624 66880 26628
rect 5796 26140 5860 26144
rect 5796 26084 5800 26140
rect 5800 26084 5856 26140
rect 5856 26084 5860 26140
rect 5796 26080 5860 26084
rect 5876 26140 5940 26144
rect 5876 26084 5880 26140
rect 5880 26084 5936 26140
rect 5936 26084 5940 26140
rect 5876 26080 5940 26084
rect 5956 26140 6020 26144
rect 5956 26084 5960 26140
rect 5960 26084 6016 26140
rect 6016 26084 6020 26140
rect 5956 26080 6020 26084
rect 6036 26140 6100 26144
rect 6036 26084 6040 26140
rect 6040 26084 6096 26140
rect 6096 26084 6100 26140
rect 6036 26080 6100 26084
rect 36516 26140 36580 26144
rect 36516 26084 36520 26140
rect 36520 26084 36576 26140
rect 36576 26084 36580 26140
rect 36516 26080 36580 26084
rect 36596 26140 36660 26144
rect 36596 26084 36600 26140
rect 36600 26084 36656 26140
rect 36656 26084 36660 26140
rect 36596 26080 36660 26084
rect 36676 26140 36740 26144
rect 36676 26084 36680 26140
rect 36680 26084 36736 26140
rect 36736 26084 36740 26140
rect 36676 26080 36740 26084
rect 36756 26140 36820 26144
rect 36756 26084 36760 26140
rect 36760 26084 36816 26140
rect 36816 26084 36820 26140
rect 36756 26080 36820 26084
rect 67236 26140 67300 26144
rect 67236 26084 67240 26140
rect 67240 26084 67296 26140
rect 67296 26084 67300 26140
rect 67236 26080 67300 26084
rect 67316 26140 67380 26144
rect 67316 26084 67320 26140
rect 67320 26084 67376 26140
rect 67376 26084 67380 26140
rect 67316 26080 67380 26084
rect 67396 26140 67460 26144
rect 67396 26084 67400 26140
rect 67400 26084 67456 26140
rect 67456 26084 67460 26140
rect 67396 26080 67460 26084
rect 67476 26140 67540 26144
rect 67476 26084 67480 26140
rect 67480 26084 67536 26140
rect 67536 26084 67540 26140
rect 67476 26080 67540 26084
rect 5136 25596 5200 25600
rect 5136 25540 5140 25596
rect 5140 25540 5196 25596
rect 5196 25540 5200 25596
rect 5136 25536 5200 25540
rect 5216 25596 5280 25600
rect 5216 25540 5220 25596
rect 5220 25540 5276 25596
rect 5276 25540 5280 25596
rect 5216 25536 5280 25540
rect 5296 25596 5360 25600
rect 5296 25540 5300 25596
rect 5300 25540 5356 25596
rect 5356 25540 5360 25596
rect 5296 25536 5360 25540
rect 5376 25596 5440 25600
rect 5376 25540 5380 25596
rect 5380 25540 5436 25596
rect 5436 25540 5440 25596
rect 5376 25536 5440 25540
rect 35856 25596 35920 25600
rect 35856 25540 35860 25596
rect 35860 25540 35916 25596
rect 35916 25540 35920 25596
rect 35856 25536 35920 25540
rect 35936 25596 36000 25600
rect 35936 25540 35940 25596
rect 35940 25540 35996 25596
rect 35996 25540 36000 25596
rect 35936 25536 36000 25540
rect 36016 25596 36080 25600
rect 36016 25540 36020 25596
rect 36020 25540 36076 25596
rect 36076 25540 36080 25596
rect 36016 25536 36080 25540
rect 36096 25596 36160 25600
rect 36096 25540 36100 25596
rect 36100 25540 36156 25596
rect 36156 25540 36160 25596
rect 36096 25536 36160 25540
rect 66576 25596 66640 25600
rect 66576 25540 66580 25596
rect 66580 25540 66636 25596
rect 66636 25540 66640 25596
rect 66576 25536 66640 25540
rect 66656 25596 66720 25600
rect 66656 25540 66660 25596
rect 66660 25540 66716 25596
rect 66716 25540 66720 25596
rect 66656 25536 66720 25540
rect 66736 25596 66800 25600
rect 66736 25540 66740 25596
rect 66740 25540 66796 25596
rect 66796 25540 66800 25596
rect 66736 25536 66800 25540
rect 66816 25596 66880 25600
rect 66816 25540 66820 25596
rect 66820 25540 66876 25596
rect 66876 25540 66880 25596
rect 66816 25536 66880 25540
rect 5796 25052 5860 25056
rect 5796 24996 5800 25052
rect 5800 24996 5856 25052
rect 5856 24996 5860 25052
rect 5796 24992 5860 24996
rect 5876 25052 5940 25056
rect 5876 24996 5880 25052
rect 5880 24996 5936 25052
rect 5936 24996 5940 25052
rect 5876 24992 5940 24996
rect 5956 25052 6020 25056
rect 5956 24996 5960 25052
rect 5960 24996 6016 25052
rect 6016 24996 6020 25052
rect 5956 24992 6020 24996
rect 6036 25052 6100 25056
rect 6036 24996 6040 25052
rect 6040 24996 6096 25052
rect 6096 24996 6100 25052
rect 6036 24992 6100 24996
rect 36516 25052 36580 25056
rect 36516 24996 36520 25052
rect 36520 24996 36576 25052
rect 36576 24996 36580 25052
rect 36516 24992 36580 24996
rect 36596 25052 36660 25056
rect 36596 24996 36600 25052
rect 36600 24996 36656 25052
rect 36656 24996 36660 25052
rect 36596 24992 36660 24996
rect 36676 25052 36740 25056
rect 36676 24996 36680 25052
rect 36680 24996 36736 25052
rect 36736 24996 36740 25052
rect 36676 24992 36740 24996
rect 36756 25052 36820 25056
rect 36756 24996 36760 25052
rect 36760 24996 36816 25052
rect 36816 24996 36820 25052
rect 36756 24992 36820 24996
rect 67236 25052 67300 25056
rect 67236 24996 67240 25052
rect 67240 24996 67296 25052
rect 67296 24996 67300 25052
rect 67236 24992 67300 24996
rect 67316 25052 67380 25056
rect 67316 24996 67320 25052
rect 67320 24996 67376 25052
rect 67376 24996 67380 25052
rect 67316 24992 67380 24996
rect 67396 25052 67460 25056
rect 67396 24996 67400 25052
rect 67400 24996 67456 25052
rect 67456 24996 67460 25052
rect 67396 24992 67460 24996
rect 67476 25052 67540 25056
rect 67476 24996 67480 25052
rect 67480 24996 67536 25052
rect 67536 24996 67540 25052
rect 67476 24992 67540 24996
rect 5136 24508 5200 24512
rect 5136 24452 5140 24508
rect 5140 24452 5196 24508
rect 5196 24452 5200 24508
rect 5136 24448 5200 24452
rect 5216 24508 5280 24512
rect 5216 24452 5220 24508
rect 5220 24452 5276 24508
rect 5276 24452 5280 24508
rect 5216 24448 5280 24452
rect 5296 24508 5360 24512
rect 5296 24452 5300 24508
rect 5300 24452 5356 24508
rect 5356 24452 5360 24508
rect 5296 24448 5360 24452
rect 5376 24508 5440 24512
rect 5376 24452 5380 24508
rect 5380 24452 5436 24508
rect 5436 24452 5440 24508
rect 5376 24448 5440 24452
rect 35856 24508 35920 24512
rect 35856 24452 35860 24508
rect 35860 24452 35916 24508
rect 35916 24452 35920 24508
rect 35856 24448 35920 24452
rect 35936 24508 36000 24512
rect 35936 24452 35940 24508
rect 35940 24452 35996 24508
rect 35996 24452 36000 24508
rect 35936 24448 36000 24452
rect 36016 24508 36080 24512
rect 36016 24452 36020 24508
rect 36020 24452 36076 24508
rect 36076 24452 36080 24508
rect 36016 24448 36080 24452
rect 36096 24508 36160 24512
rect 36096 24452 36100 24508
rect 36100 24452 36156 24508
rect 36156 24452 36160 24508
rect 36096 24448 36160 24452
rect 66576 24508 66640 24512
rect 66576 24452 66580 24508
rect 66580 24452 66636 24508
rect 66636 24452 66640 24508
rect 66576 24448 66640 24452
rect 66656 24508 66720 24512
rect 66656 24452 66660 24508
rect 66660 24452 66716 24508
rect 66716 24452 66720 24508
rect 66656 24448 66720 24452
rect 66736 24508 66800 24512
rect 66736 24452 66740 24508
rect 66740 24452 66796 24508
rect 66796 24452 66800 24508
rect 66736 24448 66800 24452
rect 66816 24508 66880 24512
rect 66816 24452 66820 24508
rect 66820 24452 66876 24508
rect 66876 24452 66880 24508
rect 66816 24448 66880 24452
rect 5796 23964 5860 23968
rect 5796 23908 5800 23964
rect 5800 23908 5856 23964
rect 5856 23908 5860 23964
rect 5796 23904 5860 23908
rect 5876 23964 5940 23968
rect 5876 23908 5880 23964
rect 5880 23908 5936 23964
rect 5936 23908 5940 23964
rect 5876 23904 5940 23908
rect 5956 23964 6020 23968
rect 5956 23908 5960 23964
rect 5960 23908 6016 23964
rect 6016 23908 6020 23964
rect 5956 23904 6020 23908
rect 6036 23964 6100 23968
rect 6036 23908 6040 23964
rect 6040 23908 6096 23964
rect 6096 23908 6100 23964
rect 6036 23904 6100 23908
rect 36516 23964 36580 23968
rect 36516 23908 36520 23964
rect 36520 23908 36576 23964
rect 36576 23908 36580 23964
rect 36516 23904 36580 23908
rect 36596 23964 36660 23968
rect 36596 23908 36600 23964
rect 36600 23908 36656 23964
rect 36656 23908 36660 23964
rect 36596 23904 36660 23908
rect 36676 23964 36740 23968
rect 36676 23908 36680 23964
rect 36680 23908 36736 23964
rect 36736 23908 36740 23964
rect 36676 23904 36740 23908
rect 36756 23964 36820 23968
rect 36756 23908 36760 23964
rect 36760 23908 36816 23964
rect 36816 23908 36820 23964
rect 36756 23904 36820 23908
rect 67236 23964 67300 23968
rect 67236 23908 67240 23964
rect 67240 23908 67296 23964
rect 67296 23908 67300 23964
rect 67236 23904 67300 23908
rect 67316 23964 67380 23968
rect 67316 23908 67320 23964
rect 67320 23908 67376 23964
rect 67376 23908 67380 23964
rect 67316 23904 67380 23908
rect 67396 23964 67460 23968
rect 67396 23908 67400 23964
rect 67400 23908 67456 23964
rect 67456 23908 67460 23964
rect 67396 23904 67460 23908
rect 67476 23964 67540 23968
rect 67476 23908 67480 23964
rect 67480 23908 67536 23964
rect 67536 23908 67540 23964
rect 67476 23904 67540 23908
rect 5136 23420 5200 23424
rect 5136 23364 5140 23420
rect 5140 23364 5196 23420
rect 5196 23364 5200 23420
rect 5136 23360 5200 23364
rect 5216 23420 5280 23424
rect 5216 23364 5220 23420
rect 5220 23364 5276 23420
rect 5276 23364 5280 23420
rect 5216 23360 5280 23364
rect 5296 23420 5360 23424
rect 5296 23364 5300 23420
rect 5300 23364 5356 23420
rect 5356 23364 5360 23420
rect 5296 23360 5360 23364
rect 5376 23420 5440 23424
rect 5376 23364 5380 23420
rect 5380 23364 5436 23420
rect 5436 23364 5440 23420
rect 5376 23360 5440 23364
rect 35856 23420 35920 23424
rect 35856 23364 35860 23420
rect 35860 23364 35916 23420
rect 35916 23364 35920 23420
rect 35856 23360 35920 23364
rect 35936 23420 36000 23424
rect 35936 23364 35940 23420
rect 35940 23364 35996 23420
rect 35996 23364 36000 23420
rect 35936 23360 36000 23364
rect 36016 23420 36080 23424
rect 36016 23364 36020 23420
rect 36020 23364 36076 23420
rect 36076 23364 36080 23420
rect 36016 23360 36080 23364
rect 36096 23420 36160 23424
rect 36096 23364 36100 23420
rect 36100 23364 36156 23420
rect 36156 23364 36160 23420
rect 36096 23360 36160 23364
rect 66576 23420 66640 23424
rect 66576 23364 66580 23420
rect 66580 23364 66636 23420
rect 66636 23364 66640 23420
rect 66576 23360 66640 23364
rect 66656 23420 66720 23424
rect 66656 23364 66660 23420
rect 66660 23364 66716 23420
rect 66716 23364 66720 23420
rect 66656 23360 66720 23364
rect 66736 23420 66800 23424
rect 66736 23364 66740 23420
rect 66740 23364 66796 23420
rect 66796 23364 66800 23420
rect 66736 23360 66800 23364
rect 66816 23420 66880 23424
rect 66816 23364 66820 23420
rect 66820 23364 66876 23420
rect 66876 23364 66880 23420
rect 66816 23360 66880 23364
rect 5796 22876 5860 22880
rect 5796 22820 5800 22876
rect 5800 22820 5856 22876
rect 5856 22820 5860 22876
rect 5796 22816 5860 22820
rect 5876 22876 5940 22880
rect 5876 22820 5880 22876
rect 5880 22820 5936 22876
rect 5936 22820 5940 22876
rect 5876 22816 5940 22820
rect 5956 22876 6020 22880
rect 5956 22820 5960 22876
rect 5960 22820 6016 22876
rect 6016 22820 6020 22876
rect 5956 22816 6020 22820
rect 6036 22876 6100 22880
rect 6036 22820 6040 22876
rect 6040 22820 6096 22876
rect 6096 22820 6100 22876
rect 6036 22816 6100 22820
rect 36516 22876 36580 22880
rect 36516 22820 36520 22876
rect 36520 22820 36576 22876
rect 36576 22820 36580 22876
rect 36516 22816 36580 22820
rect 36596 22876 36660 22880
rect 36596 22820 36600 22876
rect 36600 22820 36656 22876
rect 36656 22820 36660 22876
rect 36596 22816 36660 22820
rect 36676 22876 36740 22880
rect 36676 22820 36680 22876
rect 36680 22820 36736 22876
rect 36736 22820 36740 22876
rect 36676 22816 36740 22820
rect 36756 22876 36820 22880
rect 36756 22820 36760 22876
rect 36760 22820 36816 22876
rect 36816 22820 36820 22876
rect 36756 22816 36820 22820
rect 67236 22876 67300 22880
rect 67236 22820 67240 22876
rect 67240 22820 67296 22876
rect 67296 22820 67300 22876
rect 67236 22816 67300 22820
rect 67316 22876 67380 22880
rect 67316 22820 67320 22876
rect 67320 22820 67376 22876
rect 67376 22820 67380 22876
rect 67316 22816 67380 22820
rect 67396 22876 67460 22880
rect 67396 22820 67400 22876
rect 67400 22820 67456 22876
rect 67456 22820 67460 22876
rect 67396 22816 67460 22820
rect 67476 22876 67540 22880
rect 67476 22820 67480 22876
rect 67480 22820 67536 22876
rect 67536 22820 67540 22876
rect 67476 22816 67540 22820
rect 5136 22332 5200 22336
rect 5136 22276 5140 22332
rect 5140 22276 5196 22332
rect 5196 22276 5200 22332
rect 5136 22272 5200 22276
rect 5216 22332 5280 22336
rect 5216 22276 5220 22332
rect 5220 22276 5276 22332
rect 5276 22276 5280 22332
rect 5216 22272 5280 22276
rect 5296 22332 5360 22336
rect 5296 22276 5300 22332
rect 5300 22276 5356 22332
rect 5356 22276 5360 22332
rect 5296 22272 5360 22276
rect 5376 22332 5440 22336
rect 5376 22276 5380 22332
rect 5380 22276 5436 22332
rect 5436 22276 5440 22332
rect 5376 22272 5440 22276
rect 35856 22332 35920 22336
rect 35856 22276 35860 22332
rect 35860 22276 35916 22332
rect 35916 22276 35920 22332
rect 35856 22272 35920 22276
rect 35936 22332 36000 22336
rect 35936 22276 35940 22332
rect 35940 22276 35996 22332
rect 35996 22276 36000 22332
rect 35936 22272 36000 22276
rect 36016 22332 36080 22336
rect 36016 22276 36020 22332
rect 36020 22276 36076 22332
rect 36076 22276 36080 22332
rect 36016 22272 36080 22276
rect 36096 22332 36160 22336
rect 36096 22276 36100 22332
rect 36100 22276 36156 22332
rect 36156 22276 36160 22332
rect 36096 22272 36160 22276
rect 66576 22332 66640 22336
rect 66576 22276 66580 22332
rect 66580 22276 66636 22332
rect 66636 22276 66640 22332
rect 66576 22272 66640 22276
rect 66656 22332 66720 22336
rect 66656 22276 66660 22332
rect 66660 22276 66716 22332
rect 66716 22276 66720 22332
rect 66656 22272 66720 22276
rect 66736 22332 66800 22336
rect 66736 22276 66740 22332
rect 66740 22276 66796 22332
rect 66796 22276 66800 22332
rect 66736 22272 66800 22276
rect 66816 22332 66880 22336
rect 66816 22276 66820 22332
rect 66820 22276 66876 22332
rect 66876 22276 66880 22332
rect 66816 22272 66880 22276
rect 5796 21788 5860 21792
rect 5796 21732 5800 21788
rect 5800 21732 5856 21788
rect 5856 21732 5860 21788
rect 5796 21728 5860 21732
rect 5876 21788 5940 21792
rect 5876 21732 5880 21788
rect 5880 21732 5936 21788
rect 5936 21732 5940 21788
rect 5876 21728 5940 21732
rect 5956 21788 6020 21792
rect 5956 21732 5960 21788
rect 5960 21732 6016 21788
rect 6016 21732 6020 21788
rect 5956 21728 6020 21732
rect 6036 21788 6100 21792
rect 6036 21732 6040 21788
rect 6040 21732 6096 21788
rect 6096 21732 6100 21788
rect 6036 21728 6100 21732
rect 36516 21788 36580 21792
rect 36516 21732 36520 21788
rect 36520 21732 36576 21788
rect 36576 21732 36580 21788
rect 36516 21728 36580 21732
rect 36596 21788 36660 21792
rect 36596 21732 36600 21788
rect 36600 21732 36656 21788
rect 36656 21732 36660 21788
rect 36596 21728 36660 21732
rect 36676 21788 36740 21792
rect 36676 21732 36680 21788
rect 36680 21732 36736 21788
rect 36736 21732 36740 21788
rect 36676 21728 36740 21732
rect 36756 21788 36820 21792
rect 36756 21732 36760 21788
rect 36760 21732 36816 21788
rect 36816 21732 36820 21788
rect 36756 21728 36820 21732
rect 67236 21788 67300 21792
rect 67236 21732 67240 21788
rect 67240 21732 67296 21788
rect 67296 21732 67300 21788
rect 67236 21728 67300 21732
rect 67316 21788 67380 21792
rect 67316 21732 67320 21788
rect 67320 21732 67376 21788
rect 67376 21732 67380 21788
rect 67316 21728 67380 21732
rect 67396 21788 67460 21792
rect 67396 21732 67400 21788
rect 67400 21732 67456 21788
rect 67456 21732 67460 21788
rect 67396 21728 67460 21732
rect 67476 21788 67540 21792
rect 67476 21732 67480 21788
rect 67480 21732 67536 21788
rect 67536 21732 67540 21788
rect 67476 21728 67540 21732
rect 5136 21244 5200 21248
rect 5136 21188 5140 21244
rect 5140 21188 5196 21244
rect 5196 21188 5200 21244
rect 5136 21184 5200 21188
rect 5216 21244 5280 21248
rect 5216 21188 5220 21244
rect 5220 21188 5276 21244
rect 5276 21188 5280 21244
rect 5216 21184 5280 21188
rect 5296 21244 5360 21248
rect 5296 21188 5300 21244
rect 5300 21188 5356 21244
rect 5356 21188 5360 21244
rect 5296 21184 5360 21188
rect 5376 21244 5440 21248
rect 5376 21188 5380 21244
rect 5380 21188 5436 21244
rect 5436 21188 5440 21244
rect 5376 21184 5440 21188
rect 35856 21244 35920 21248
rect 35856 21188 35860 21244
rect 35860 21188 35916 21244
rect 35916 21188 35920 21244
rect 35856 21184 35920 21188
rect 35936 21244 36000 21248
rect 35936 21188 35940 21244
rect 35940 21188 35996 21244
rect 35996 21188 36000 21244
rect 35936 21184 36000 21188
rect 36016 21244 36080 21248
rect 36016 21188 36020 21244
rect 36020 21188 36076 21244
rect 36076 21188 36080 21244
rect 36016 21184 36080 21188
rect 36096 21244 36160 21248
rect 36096 21188 36100 21244
rect 36100 21188 36156 21244
rect 36156 21188 36160 21244
rect 36096 21184 36160 21188
rect 66576 21244 66640 21248
rect 66576 21188 66580 21244
rect 66580 21188 66636 21244
rect 66636 21188 66640 21244
rect 66576 21184 66640 21188
rect 66656 21244 66720 21248
rect 66656 21188 66660 21244
rect 66660 21188 66716 21244
rect 66716 21188 66720 21244
rect 66656 21184 66720 21188
rect 66736 21244 66800 21248
rect 66736 21188 66740 21244
rect 66740 21188 66796 21244
rect 66796 21188 66800 21244
rect 66736 21184 66800 21188
rect 66816 21244 66880 21248
rect 66816 21188 66820 21244
rect 66820 21188 66876 21244
rect 66876 21188 66880 21244
rect 66816 21184 66880 21188
rect 5796 20700 5860 20704
rect 5796 20644 5800 20700
rect 5800 20644 5856 20700
rect 5856 20644 5860 20700
rect 5796 20640 5860 20644
rect 5876 20700 5940 20704
rect 5876 20644 5880 20700
rect 5880 20644 5936 20700
rect 5936 20644 5940 20700
rect 5876 20640 5940 20644
rect 5956 20700 6020 20704
rect 5956 20644 5960 20700
rect 5960 20644 6016 20700
rect 6016 20644 6020 20700
rect 5956 20640 6020 20644
rect 6036 20700 6100 20704
rect 6036 20644 6040 20700
rect 6040 20644 6096 20700
rect 6096 20644 6100 20700
rect 6036 20640 6100 20644
rect 36516 20700 36580 20704
rect 36516 20644 36520 20700
rect 36520 20644 36576 20700
rect 36576 20644 36580 20700
rect 36516 20640 36580 20644
rect 36596 20700 36660 20704
rect 36596 20644 36600 20700
rect 36600 20644 36656 20700
rect 36656 20644 36660 20700
rect 36596 20640 36660 20644
rect 36676 20700 36740 20704
rect 36676 20644 36680 20700
rect 36680 20644 36736 20700
rect 36736 20644 36740 20700
rect 36676 20640 36740 20644
rect 36756 20700 36820 20704
rect 36756 20644 36760 20700
rect 36760 20644 36816 20700
rect 36816 20644 36820 20700
rect 36756 20640 36820 20644
rect 67236 20700 67300 20704
rect 67236 20644 67240 20700
rect 67240 20644 67296 20700
rect 67296 20644 67300 20700
rect 67236 20640 67300 20644
rect 67316 20700 67380 20704
rect 67316 20644 67320 20700
rect 67320 20644 67376 20700
rect 67376 20644 67380 20700
rect 67316 20640 67380 20644
rect 67396 20700 67460 20704
rect 67396 20644 67400 20700
rect 67400 20644 67456 20700
rect 67456 20644 67460 20700
rect 67396 20640 67460 20644
rect 67476 20700 67540 20704
rect 67476 20644 67480 20700
rect 67480 20644 67536 20700
rect 67536 20644 67540 20700
rect 67476 20640 67540 20644
rect 5136 20156 5200 20160
rect 5136 20100 5140 20156
rect 5140 20100 5196 20156
rect 5196 20100 5200 20156
rect 5136 20096 5200 20100
rect 5216 20156 5280 20160
rect 5216 20100 5220 20156
rect 5220 20100 5276 20156
rect 5276 20100 5280 20156
rect 5216 20096 5280 20100
rect 5296 20156 5360 20160
rect 5296 20100 5300 20156
rect 5300 20100 5356 20156
rect 5356 20100 5360 20156
rect 5296 20096 5360 20100
rect 5376 20156 5440 20160
rect 5376 20100 5380 20156
rect 5380 20100 5436 20156
rect 5436 20100 5440 20156
rect 5376 20096 5440 20100
rect 35856 20156 35920 20160
rect 35856 20100 35860 20156
rect 35860 20100 35916 20156
rect 35916 20100 35920 20156
rect 35856 20096 35920 20100
rect 35936 20156 36000 20160
rect 35936 20100 35940 20156
rect 35940 20100 35996 20156
rect 35996 20100 36000 20156
rect 35936 20096 36000 20100
rect 36016 20156 36080 20160
rect 36016 20100 36020 20156
rect 36020 20100 36076 20156
rect 36076 20100 36080 20156
rect 36016 20096 36080 20100
rect 36096 20156 36160 20160
rect 36096 20100 36100 20156
rect 36100 20100 36156 20156
rect 36156 20100 36160 20156
rect 36096 20096 36160 20100
rect 66576 20156 66640 20160
rect 66576 20100 66580 20156
rect 66580 20100 66636 20156
rect 66636 20100 66640 20156
rect 66576 20096 66640 20100
rect 66656 20156 66720 20160
rect 66656 20100 66660 20156
rect 66660 20100 66716 20156
rect 66716 20100 66720 20156
rect 66656 20096 66720 20100
rect 66736 20156 66800 20160
rect 66736 20100 66740 20156
rect 66740 20100 66796 20156
rect 66796 20100 66800 20156
rect 66736 20096 66800 20100
rect 66816 20156 66880 20160
rect 66816 20100 66820 20156
rect 66820 20100 66876 20156
rect 66876 20100 66880 20156
rect 66816 20096 66880 20100
rect 5796 19612 5860 19616
rect 5796 19556 5800 19612
rect 5800 19556 5856 19612
rect 5856 19556 5860 19612
rect 5796 19552 5860 19556
rect 5876 19612 5940 19616
rect 5876 19556 5880 19612
rect 5880 19556 5936 19612
rect 5936 19556 5940 19612
rect 5876 19552 5940 19556
rect 5956 19612 6020 19616
rect 5956 19556 5960 19612
rect 5960 19556 6016 19612
rect 6016 19556 6020 19612
rect 5956 19552 6020 19556
rect 6036 19612 6100 19616
rect 6036 19556 6040 19612
rect 6040 19556 6096 19612
rect 6096 19556 6100 19612
rect 6036 19552 6100 19556
rect 36516 19612 36580 19616
rect 36516 19556 36520 19612
rect 36520 19556 36576 19612
rect 36576 19556 36580 19612
rect 36516 19552 36580 19556
rect 36596 19612 36660 19616
rect 36596 19556 36600 19612
rect 36600 19556 36656 19612
rect 36656 19556 36660 19612
rect 36596 19552 36660 19556
rect 36676 19612 36740 19616
rect 36676 19556 36680 19612
rect 36680 19556 36736 19612
rect 36736 19556 36740 19612
rect 36676 19552 36740 19556
rect 36756 19612 36820 19616
rect 36756 19556 36760 19612
rect 36760 19556 36816 19612
rect 36816 19556 36820 19612
rect 36756 19552 36820 19556
rect 67236 19612 67300 19616
rect 67236 19556 67240 19612
rect 67240 19556 67296 19612
rect 67296 19556 67300 19612
rect 67236 19552 67300 19556
rect 67316 19612 67380 19616
rect 67316 19556 67320 19612
rect 67320 19556 67376 19612
rect 67376 19556 67380 19612
rect 67316 19552 67380 19556
rect 67396 19612 67460 19616
rect 67396 19556 67400 19612
rect 67400 19556 67456 19612
rect 67456 19556 67460 19612
rect 67396 19552 67460 19556
rect 67476 19612 67540 19616
rect 67476 19556 67480 19612
rect 67480 19556 67536 19612
rect 67536 19556 67540 19612
rect 67476 19552 67540 19556
rect 5136 19068 5200 19072
rect 5136 19012 5140 19068
rect 5140 19012 5196 19068
rect 5196 19012 5200 19068
rect 5136 19008 5200 19012
rect 5216 19068 5280 19072
rect 5216 19012 5220 19068
rect 5220 19012 5276 19068
rect 5276 19012 5280 19068
rect 5216 19008 5280 19012
rect 5296 19068 5360 19072
rect 5296 19012 5300 19068
rect 5300 19012 5356 19068
rect 5356 19012 5360 19068
rect 5296 19008 5360 19012
rect 5376 19068 5440 19072
rect 5376 19012 5380 19068
rect 5380 19012 5436 19068
rect 5436 19012 5440 19068
rect 5376 19008 5440 19012
rect 35856 19068 35920 19072
rect 35856 19012 35860 19068
rect 35860 19012 35916 19068
rect 35916 19012 35920 19068
rect 35856 19008 35920 19012
rect 35936 19068 36000 19072
rect 35936 19012 35940 19068
rect 35940 19012 35996 19068
rect 35996 19012 36000 19068
rect 35936 19008 36000 19012
rect 36016 19068 36080 19072
rect 36016 19012 36020 19068
rect 36020 19012 36076 19068
rect 36076 19012 36080 19068
rect 36016 19008 36080 19012
rect 36096 19068 36160 19072
rect 36096 19012 36100 19068
rect 36100 19012 36156 19068
rect 36156 19012 36160 19068
rect 36096 19008 36160 19012
rect 66576 19068 66640 19072
rect 66576 19012 66580 19068
rect 66580 19012 66636 19068
rect 66636 19012 66640 19068
rect 66576 19008 66640 19012
rect 66656 19068 66720 19072
rect 66656 19012 66660 19068
rect 66660 19012 66716 19068
rect 66716 19012 66720 19068
rect 66656 19008 66720 19012
rect 66736 19068 66800 19072
rect 66736 19012 66740 19068
rect 66740 19012 66796 19068
rect 66796 19012 66800 19068
rect 66736 19008 66800 19012
rect 66816 19068 66880 19072
rect 66816 19012 66820 19068
rect 66820 19012 66876 19068
rect 66876 19012 66880 19068
rect 66816 19008 66880 19012
rect 5796 18524 5860 18528
rect 5796 18468 5800 18524
rect 5800 18468 5856 18524
rect 5856 18468 5860 18524
rect 5796 18464 5860 18468
rect 5876 18524 5940 18528
rect 5876 18468 5880 18524
rect 5880 18468 5936 18524
rect 5936 18468 5940 18524
rect 5876 18464 5940 18468
rect 5956 18524 6020 18528
rect 5956 18468 5960 18524
rect 5960 18468 6016 18524
rect 6016 18468 6020 18524
rect 5956 18464 6020 18468
rect 6036 18524 6100 18528
rect 6036 18468 6040 18524
rect 6040 18468 6096 18524
rect 6096 18468 6100 18524
rect 6036 18464 6100 18468
rect 36516 18524 36580 18528
rect 36516 18468 36520 18524
rect 36520 18468 36576 18524
rect 36576 18468 36580 18524
rect 36516 18464 36580 18468
rect 36596 18524 36660 18528
rect 36596 18468 36600 18524
rect 36600 18468 36656 18524
rect 36656 18468 36660 18524
rect 36596 18464 36660 18468
rect 36676 18524 36740 18528
rect 36676 18468 36680 18524
rect 36680 18468 36736 18524
rect 36736 18468 36740 18524
rect 36676 18464 36740 18468
rect 36756 18524 36820 18528
rect 36756 18468 36760 18524
rect 36760 18468 36816 18524
rect 36816 18468 36820 18524
rect 36756 18464 36820 18468
rect 67236 18524 67300 18528
rect 67236 18468 67240 18524
rect 67240 18468 67296 18524
rect 67296 18468 67300 18524
rect 67236 18464 67300 18468
rect 67316 18524 67380 18528
rect 67316 18468 67320 18524
rect 67320 18468 67376 18524
rect 67376 18468 67380 18524
rect 67316 18464 67380 18468
rect 67396 18524 67460 18528
rect 67396 18468 67400 18524
rect 67400 18468 67456 18524
rect 67456 18468 67460 18524
rect 67396 18464 67460 18468
rect 67476 18524 67540 18528
rect 67476 18468 67480 18524
rect 67480 18468 67536 18524
rect 67536 18468 67540 18524
rect 67476 18464 67540 18468
rect 5136 17980 5200 17984
rect 5136 17924 5140 17980
rect 5140 17924 5196 17980
rect 5196 17924 5200 17980
rect 5136 17920 5200 17924
rect 5216 17980 5280 17984
rect 5216 17924 5220 17980
rect 5220 17924 5276 17980
rect 5276 17924 5280 17980
rect 5216 17920 5280 17924
rect 5296 17980 5360 17984
rect 5296 17924 5300 17980
rect 5300 17924 5356 17980
rect 5356 17924 5360 17980
rect 5296 17920 5360 17924
rect 5376 17980 5440 17984
rect 5376 17924 5380 17980
rect 5380 17924 5436 17980
rect 5436 17924 5440 17980
rect 5376 17920 5440 17924
rect 35856 17980 35920 17984
rect 35856 17924 35860 17980
rect 35860 17924 35916 17980
rect 35916 17924 35920 17980
rect 35856 17920 35920 17924
rect 35936 17980 36000 17984
rect 35936 17924 35940 17980
rect 35940 17924 35996 17980
rect 35996 17924 36000 17980
rect 35936 17920 36000 17924
rect 36016 17980 36080 17984
rect 36016 17924 36020 17980
rect 36020 17924 36076 17980
rect 36076 17924 36080 17980
rect 36016 17920 36080 17924
rect 36096 17980 36160 17984
rect 36096 17924 36100 17980
rect 36100 17924 36156 17980
rect 36156 17924 36160 17980
rect 36096 17920 36160 17924
rect 66576 17980 66640 17984
rect 66576 17924 66580 17980
rect 66580 17924 66636 17980
rect 66636 17924 66640 17980
rect 66576 17920 66640 17924
rect 66656 17980 66720 17984
rect 66656 17924 66660 17980
rect 66660 17924 66716 17980
rect 66716 17924 66720 17980
rect 66656 17920 66720 17924
rect 66736 17980 66800 17984
rect 66736 17924 66740 17980
rect 66740 17924 66796 17980
rect 66796 17924 66800 17980
rect 66736 17920 66800 17924
rect 66816 17980 66880 17984
rect 66816 17924 66820 17980
rect 66820 17924 66876 17980
rect 66876 17924 66880 17980
rect 66816 17920 66880 17924
rect 5796 17436 5860 17440
rect 5796 17380 5800 17436
rect 5800 17380 5856 17436
rect 5856 17380 5860 17436
rect 5796 17376 5860 17380
rect 5876 17436 5940 17440
rect 5876 17380 5880 17436
rect 5880 17380 5936 17436
rect 5936 17380 5940 17436
rect 5876 17376 5940 17380
rect 5956 17436 6020 17440
rect 5956 17380 5960 17436
rect 5960 17380 6016 17436
rect 6016 17380 6020 17436
rect 5956 17376 6020 17380
rect 6036 17436 6100 17440
rect 6036 17380 6040 17436
rect 6040 17380 6096 17436
rect 6096 17380 6100 17436
rect 6036 17376 6100 17380
rect 36516 17436 36580 17440
rect 36516 17380 36520 17436
rect 36520 17380 36576 17436
rect 36576 17380 36580 17436
rect 36516 17376 36580 17380
rect 36596 17436 36660 17440
rect 36596 17380 36600 17436
rect 36600 17380 36656 17436
rect 36656 17380 36660 17436
rect 36596 17376 36660 17380
rect 36676 17436 36740 17440
rect 36676 17380 36680 17436
rect 36680 17380 36736 17436
rect 36736 17380 36740 17436
rect 36676 17376 36740 17380
rect 36756 17436 36820 17440
rect 36756 17380 36760 17436
rect 36760 17380 36816 17436
rect 36816 17380 36820 17436
rect 36756 17376 36820 17380
rect 67236 17436 67300 17440
rect 67236 17380 67240 17436
rect 67240 17380 67296 17436
rect 67296 17380 67300 17436
rect 67236 17376 67300 17380
rect 67316 17436 67380 17440
rect 67316 17380 67320 17436
rect 67320 17380 67376 17436
rect 67376 17380 67380 17436
rect 67316 17376 67380 17380
rect 67396 17436 67460 17440
rect 67396 17380 67400 17436
rect 67400 17380 67456 17436
rect 67456 17380 67460 17436
rect 67396 17376 67460 17380
rect 67476 17436 67540 17440
rect 67476 17380 67480 17436
rect 67480 17380 67536 17436
rect 67536 17380 67540 17436
rect 67476 17376 67540 17380
rect 5136 16892 5200 16896
rect 5136 16836 5140 16892
rect 5140 16836 5196 16892
rect 5196 16836 5200 16892
rect 5136 16832 5200 16836
rect 5216 16892 5280 16896
rect 5216 16836 5220 16892
rect 5220 16836 5276 16892
rect 5276 16836 5280 16892
rect 5216 16832 5280 16836
rect 5296 16892 5360 16896
rect 5296 16836 5300 16892
rect 5300 16836 5356 16892
rect 5356 16836 5360 16892
rect 5296 16832 5360 16836
rect 5376 16892 5440 16896
rect 5376 16836 5380 16892
rect 5380 16836 5436 16892
rect 5436 16836 5440 16892
rect 5376 16832 5440 16836
rect 35856 16892 35920 16896
rect 35856 16836 35860 16892
rect 35860 16836 35916 16892
rect 35916 16836 35920 16892
rect 35856 16832 35920 16836
rect 35936 16892 36000 16896
rect 35936 16836 35940 16892
rect 35940 16836 35996 16892
rect 35996 16836 36000 16892
rect 35936 16832 36000 16836
rect 36016 16892 36080 16896
rect 36016 16836 36020 16892
rect 36020 16836 36076 16892
rect 36076 16836 36080 16892
rect 36016 16832 36080 16836
rect 36096 16892 36160 16896
rect 36096 16836 36100 16892
rect 36100 16836 36156 16892
rect 36156 16836 36160 16892
rect 36096 16832 36160 16836
rect 66576 16892 66640 16896
rect 66576 16836 66580 16892
rect 66580 16836 66636 16892
rect 66636 16836 66640 16892
rect 66576 16832 66640 16836
rect 66656 16892 66720 16896
rect 66656 16836 66660 16892
rect 66660 16836 66716 16892
rect 66716 16836 66720 16892
rect 66656 16832 66720 16836
rect 66736 16892 66800 16896
rect 66736 16836 66740 16892
rect 66740 16836 66796 16892
rect 66796 16836 66800 16892
rect 66736 16832 66800 16836
rect 66816 16892 66880 16896
rect 66816 16836 66820 16892
rect 66820 16836 66876 16892
rect 66876 16836 66880 16892
rect 66816 16832 66880 16836
rect 5796 16348 5860 16352
rect 5796 16292 5800 16348
rect 5800 16292 5856 16348
rect 5856 16292 5860 16348
rect 5796 16288 5860 16292
rect 5876 16348 5940 16352
rect 5876 16292 5880 16348
rect 5880 16292 5936 16348
rect 5936 16292 5940 16348
rect 5876 16288 5940 16292
rect 5956 16348 6020 16352
rect 5956 16292 5960 16348
rect 5960 16292 6016 16348
rect 6016 16292 6020 16348
rect 5956 16288 6020 16292
rect 6036 16348 6100 16352
rect 6036 16292 6040 16348
rect 6040 16292 6096 16348
rect 6096 16292 6100 16348
rect 6036 16288 6100 16292
rect 36516 16348 36580 16352
rect 36516 16292 36520 16348
rect 36520 16292 36576 16348
rect 36576 16292 36580 16348
rect 36516 16288 36580 16292
rect 36596 16348 36660 16352
rect 36596 16292 36600 16348
rect 36600 16292 36656 16348
rect 36656 16292 36660 16348
rect 36596 16288 36660 16292
rect 36676 16348 36740 16352
rect 36676 16292 36680 16348
rect 36680 16292 36736 16348
rect 36736 16292 36740 16348
rect 36676 16288 36740 16292
rect 36756 16348 36820 16352
rect 36756 16292 36760 16348
rect 36760 16292 36816 16348
rect 36816 16292 36820 16348
rect 36756 16288 36820 16292
rect 67236 16348 67300 16352
rect 67236 16292 67240 16348
rect 67240 16292 67296 16348
rect 67296 16292 67300 16348
rect 67236 16288 67300 16292
rect 67316 16348 67380 16352
rect 67316 16292 67320 16348
rect 67320 16292 67376 16348
rect 67376 16292 67380 16348
rect 67316 16288 67380 16292
rect 67396 16348 67460 16352
rect 67396 16292 67400 16348
rect 67400 16292 67456 16348
rect 67456 16292 67460 16348
rect 67396 16288 67460 16292
rect 67476 16348 67540 16352
rect 67476 16292 67480 16348
rect 67480 16292 67536 16348
rect 67536 16292 67540 16348
rect 67476 16288 67540 16292
rect 5136 15804 5200 15808
rect 5136 15748 5140 15804
rect 5140 15748 5196 15804
rect 5196 15748 5200 15804
rect 5136 15744 5200 15748
rect 5216 15804 5280 15808
rect 5216 15748 5220 15804
rect 5220 15748 5276 15804
rect 5276 15748 5280 15804
rect 5216 15744 5280 15748
rect 5296 15804 5360 15808
rect 5296 15748 5300 15804
rect 5300 15748 5356 15804
rect 5356 15748 5360 15804
rect 5296 15744 5360 15748
rect 5376 15804 5440 15808
rect 5376 15748 5380 15804
rect 5380 15748 5436 15804
rect 5436 15748 5440 15804
rect 5376 15744 5440 15748
rect 35856 15804 35920 15808
rect 35856 15748 35860 15804
rect 35860 15748 35916 15804
rect 35916 15748 35920 15804
rect 35856 15744 35920 15748
rect 35936 15804 36000 15808
rect 35936 15748 35940 15804
rect 35940 15748 35996 15804
rect 35996 15748 36000 15804
rect 35936 15744 36000 15748
rect 36016 15804 36080 15808
rect 36016 15748 36020 15804
rect 36020 15748 36076 15804
rect 36076 15748 36080 15804
rect 36016 15744 36080 15748
rect 36096 15804 36160 15808
rect 36096 15748 36100 15804
rect 36100 15748 36156 15804
rect 36156 15748 36160 15804
rect 36096 15744 36160 15748
rect 66576 15804 66640 15808
rect 66576 15748 66580 15804
rect 66580 15748 66636 15804
rect 66636 15748 66640 15804
rect 66576 15744 66640 15748
rect 66656 15804 66720 15808
rect 66656 15748 66660 15804
rect 66660 15748 66716 15804
rect 66716 15748 66720 15804
rect 66656 15744 66720 15748
rect 66736 15804 66800 15808
rect 66736 15748 66740 15804
rect 66740 15748 66796 15804
rect 66796 15748 66800 15804
rect 66736 15744 66800 15748
rect 66816 15804 66880 15808
rect 66816 15748 66820 15804
rect 66820 15748 66876 15804
rect 66876 15748 66880 15804
rect 66816 15744 66880 15748
rect 5796 15260 5860 15264
rect 5796 15204 5800 15260
rect 5800 15204 5856 15260
rect 5856 15204 5860 15260
rect 5796 15200 5860 15204
rect 5876 15260 5940 15264
rect 5876 15204 5880 15260
rect 5880 15204 5936 15260
rect 5936 15204 5940 15260
rect 5876 15200 5940 15204
rect 5956 15260 6020 15264
rect 5956 15204 5960 15260
rect 5960 15204 6016 15260
rect 6016 15204 6020 15260
rect 5956 15200 6020 15204
rect 6036 15260 6100 15264
rect 6036 15204 6040 15260
rect 6040 15204 6096 15260
rect 6096 15204 6100 15260
rect 6036 15200 6100 15204
rect 36516 15260 36580 15264
rect 36516 15204 36520 15260
rect 36520 15204 36576 15260
rect 36576 15204 36580 15260
rect 36516 15200 36580 15204
rect 36596 15260 36660 15264
rect 36596 15204 36600 15260
rect 36600 15204 36656 15260
rect 36656 15204 36660 15260
rect 36596 15200 36660 15204
rect 36676 15260 36740 15264
rect 36676 15204 36680 15260
rect 36680 15204 36736 15260
rect 36736 15204 36740 15260
rect 36676 15200 36740 15204
rect 36756 15260 36820 15264
rect 36756 15204 36760 15260
rect 36760 15204 36816 15260
rect 36816 15204 36820 15260
rect 36756 15200 36820 15204
rect 67236 15260 67300 15264
rect 67236 15204 67240 15260
rect 67240 15204 67296 15260
rect 67296 15204 67300 15260
rect 67236 15200 67300 15204
rect 67316 15260 67380 15264
rect 67316 15204 67320 15260
rect 67320 15204 67376 15260
rect 67376 15204 67380 15260
rect 67316 15200 67380 15204
rect 67396 15260 67460 15264
rect 67396 15204 67400 15260
rect 67400 15204 67456 15260
rect 67456 15204 67460 15260
rect 67396 15200 67460 15204
rect 67476 15260 67540 15264
rect 67476 15204 67480 15260
rect 67480 15204 67536 15260
rect 67536 15204 67540 15260
rect 67476 15200 67540 15204
rect 5136 14716 5200 14720
rect 5136 14660 5140 14716
rect 5140 14660 5196 14716
rect 5196 14660 5200 14716
rect 5136 14656 5200 14660
rect 5216 14716 5280 14720
rect 5216 14660 5220 14716
rect 5220 14660 5276 14716
rect 5276 14660 5280 14716
rect 5216 14656 5280 14660
rect 5296 14716 5360 14720
rect 5296 14660 5300 14716
rect 5300 14660 5356 14716
rect 5356 14660 5360 14716
rect 5296 14656 5360 14660
rect 5376 14716 5440 14720
rect 5376 14660 5380 14716
rect 5380 14660 5436 14716
rect 5436 14660 5440 14716
rect 5376 14656 5440 14660
rect 35856 14716 35920 14720
rect 35856 14660 35860 14716
rect 35860 14660 35916 14716
rect 35916 14660 35920 14716
rect 35856 14656 35920 14660
rect 35936 14716 36000 14720
rect 35936 14660 35940 14716
rect 35940 14660 35996 14716
rect 35996 14660 36000 14716
rect 35936 14656 36000 14660
rect 36016 14716 36080 14720
rect 36016 14660 36020 14716
rect 36020 14660 36076 14716
rect 36076 14660 36080 14716
rect 36016 14656 36080 14660
rect 36096 14716 36160 14720
rect 36096 14660 36100 14716
rect 36100 14660 36156 14716
rect 36156 14660 36160 14716
rect 36096 14656 36160 14660
rect 66576 14716 66640 14720
rect 66576 14660 66580 14716
rect 66580 14660 66636 14716
rect 66636 14660 66640 14716
rect 66576 14656 66640 14660
rect 66656 14716 66720 14720
rect 66656 14660 66660 14716
rect 66660 14660 66716 14716
rect 66716 14660 66720 14716
rect 66656 14656 66720 14660
rect 66736 14716 66800 14720
rect 66736 14660 66740 14716
rect 66740 14660 66796 14716
rect 66796 14660 66800 14716
rect 66736 14656 66800 14660
rect 66816 14716 66880 14720
rect 66816 14660 66820 14716
rect 66820 14660 66876 14716
rect 66876 14660 66880 14716
rect 66816 14656 66880 14660
rect 5796 14172 5860 14176
rect 5796 14116 5800 14172
rect 5800 14116 5856 14172
rect 5856 14116 5860 14172
rect 5796 14112 5860 14116
rect 5876 14172 5940 14176
rect 5876 14116 5880 14172
rect 5880 14116 5936 14172
rect 5936 14116 5940 14172
rect 5876 14112 5940 14116
rect 5956 14172 6020 14176
rect 5956 14116 5960 14172
rect 5960 14116 6016 14172
rect 6016 14116 6020 14172
rect 5956 14112 6020 14116
rect 6036 14172 6100 14176
rect 6036 14116 6040 14172
rect 6040 14116 6096 14172
rect 6096 14116 6100 14172
rect 6036 14112 6100 14116
rect 36516 14172 36580 14176
rect 36516 14116 36520 14172
rect 36520 14116 36576 14172
rect 36576 14116 36580 14172
rect 36516 14112 36580 14116
rect 36596 14172 36660 14176
rect 36596 14116 36600 14172
rect 36600 14116 36656 14172
rect 36656 14116 36660 14172
rect 36596 14112 36660 14116
rect 36676 14172 36740 14176
rect 36676 14116 36680 14172
rect 36680 14116 36736 14172
rect 36736 14116 36740 14172
rect 36676 14112 36740 14116
rect 36756 14172 36820 14176
rect 36756 14116 36760 14172
rect 36760 14116 36816 14172
rect 36816 14116 36820 14172
rect 36756 14112 36820 14116
rect 67236 14172 67300 14176
rect 67236 14116 67240 14172
rect 67240 14116 67296 14172
rect 67296 14116 67300 14172
rect 67236 14112 67300 14116
rect 67316 14172 67380 14176
rect 67316 14116 67320 14172
rect 67320 14116 67376 14172
rect 67376 14116 67380 14172
rect 67316 14112 67380 14116
rect 67396 14172 67460 14176
rect 67396 14116 67400 14172
rect 67400 14116 67456 14172
rect 67456 14116 67460 14172
rect 67396 14112 67460 14116
rect 67476 14172 67540 14176
rect 67476 14116 67480 14172
rect 67480 14116 67536 14172
rect 67536 14116 67540 14172
rect 67476 14112 67540 14116
rect 5136 13628 5200 13632
rect 5136 13572 5140 13628
rect 5140 13572 5196 13628
rect 5196 13572 5200 13628
rect 5136 13568 5200 13572
rect 5216 13628 5280 13632
rect 5216 13572 5220 13628
rect 5220 13572 5276 13628
rect 5276 13572 5280 13628
rect 5216 13568 5280 13572
rect 5296 13628 5360 13632
rect 5296 13572 5300 13628
rect 5300 13572 5356 13628
rect 5356 13572 5360 13628
rect 5296 13568 5360 13572
rect 5376 13628 5440 13632
rect 5376 13572 5380 13628
rect 5380 13572 5436 13628
rect 5436 13572 5440 13628
rect 5376 13568 5440 13572
rect 35856 13628 35920 13632
rect 35856 13572 35860 13628
rect 35860 13572 35916 13628
rect 35916 13572 35920 13628
rect 35856 13568 35920 13572
rect 35936 13628 36000 13632
rect 35936 13572 35940 13628
rect 35940 13572 35996 13628
rect 35996 13572 36000 13628
rect 35936 13568 36000 13572
rect 36016 13628 36080 13632
rect 36016 13572 36020 13628
rect 36020 13572 36076 13628
rect 36076 13572 36080 13628
rect 36016 13568 36080 13572
rect 36096 13628 36160 13632
rect 36096 13572 36100 13628
rect 36100 13572 36156 13628
rect 36156 13572 36160 13628
rect 36096 13568 36160 13572
rect 66576 13628 66640 13632
rect 66576 13572 66580 13628
rect 66580 13572 66636 13628
rect 66636 13572 66640 13628
rect 66576 13568 66640 13572
rect 66656 13628 66720 13632
rect 66656 13572 66660 13628
rect 66660 13572 66716 13628
rect 66716 13572 66720 13628
rect 66656 13568 66720 13572
rect 66736 13628 66800 13632
rect 66736 13572 66740 13628
rect 66740 13572 66796 13628
rect 66796 13572 66800 13628
rect 66736 13568 66800 13572
rect 66816 13628 66880 13632
rect 66816 13572 66820 13628
rect 66820 13572 66876 13628
rect 66876 13572 66880 13628
rect 66816 13568 66880 13572
rect 5796 13084 5860 13088
rect 5796 13028 5800 13084
rect 5800 13028 5856 13084
rect 5856 13028 5860 13084
rect 5796 13024 5860 13028
rect 5876 13084 5940 13088
rect 5876 13028 5880 13084
rect 5880 13028 5936 13084
rect 5936 13028 5940 13084
rect 5876 13024 5940 13028
rect 5956 13084 6020 13088
rect 5956 13028 5960 13084
rect 5960 13028 6016 13084
rect 6016 13028 6020 13084
rect 5956 13024 6020 13028
rect 6036 13084 6100 13088
rect 6036 13028 6040 13084
rect 6040 13028 6096 13084
rect 6096 13028 6100 13084
rect 6036 13024 6100 13028
rect 36516 13084 36580 13088
rect 36516 13028 36520 13084
rect 36520 13028 36576 13084
rect 36576 13028 36580 13084
rect 36516 13024 36580 13028
rect 36596 13084 36660 13088
rect 36596 13028 36600 13084
rect 36600 13028 36656 13084
rect 36656 13028 36660 13084
rect 36596 13024 36660 13028
rect 36676 13084 36740 13088
rect 36676 13028 36680 13084
rect 36680 13028 36736 13084
rect 36736 13028 36740 13084
rect 36676 13024 36740 13028
rect 36756 13084 36820 13088
rect 36756 13028 36760 13084
rect 36760 13028 36816 13084
rect 36816 13028 36820 13084
rect 36756 13024 36820 13028
rect 67236 13084 67300 13088
rect 67236 13028 67240 13084
rect 67240 13028 67296 13084
rect 67296 13028 67300 13084
rect 67236 13024 67300 13028
rect 67316 13084 67380 13088
rect 67316 13028 67320 13084
rect 67320 13028 67376 13084
rect 67376 13028 67380 13084
rect 67316 13024 67380 13028
rect 67396 13084 67460 13088
rect 67396 13028 67400 13084
rect 67400 13028 67456 13084
rect 67456 13028 67460 13084
rect 67396 13024 67460 13028
rect 67476 13084 67540 13088
rect 67476 13028 67480 13084
rect 67480 13028 67536 13084
rect 67536 13028 67540 13084
rect 67476 13024 67540 13028
rect 5136 12540 5200 12544
rect 5136 12484 5140 12540
rect 5140 12484 5196 12540
rect 5196 12484 5200 12540
rect 5136 12480 5200 12484
rect 5216 12540 5280 12544
rect 5216 12484 5220 12540
rect 5220 12484 5276 12540
rect 5276 12484 5280 12540
rect 5216 12480 5280 12484
rect 5296 12540 5360 12544
rect 5296 12484 5300 12540
rect 5300 12484 5356 12540
rect 5356 12484 5360 12540
rect 5296 12480 5360 12484
rect 5376 12540 5440 12544
rect 5376 12484 5380 12540
rect 5380 12484 5436 12540
rect 5436 12484 5440 12540
rect 5376 12480 5440 12484
rect 35856 12540 35920 12544
rect 35856 12484 35860 12540
rect 35860 12484 35916 12540
rect 35916 12484 35920 12540
rect 35856 12480 35920 12484
rect 35936 12540 36000 12544
rect 35936 12484 35940 12540
rect 35940 12484 35996 12540
rect 35996 12484 36000 12540
rect 35936 12480 36000 12484
rect 36016 12540 36080 12544
rect 36016 12484 36020 12540
rect 36020 12484 36076 12540
rect 36076 12484 36080 12540
rect 36016 12480 36080 12484
rect 36096 12540 36160 12544
rect 36096 12484 36100 12540
rect 36100 12484 36156 12540
rect 36156 12484 36160 12540
rect 36096 12480 36160 12484
rect 66576 12540 66640 12544
rect 66576 12484 66580 12540
rect 66580 12484 66636 12540
rect 66636 12484 66640 12540
rect 66576 12480 66640 12484
rect 66656 12540 66720 12544
rect 66656 12484 66660 12540
rect 66660 12484 66716 12540
rect 66716 12484 66720 12540
rect 66656 12480 66720 12484
rect 66736 12540 66800 12544
rect 66736 12484 66740 12540
rect 66740 12484 66796 12540
rect 66796 12484 66800 12540
rect 66736 12480 66800 12484
rect 66816 12540 66880 12544
rect 66816 12484 66820 12540
rect 66820 12484 66876 12540
rect 66876 12484 66880 12540
rect 66816 12480 66880 12484
rect 5796 11996 5860 12000
rect 5796 11940 5800 11996
rect 5800 11940 5856 11996
rect 5856 11940 5860 11996
rect 5796 11936 5860 11940
rect 5876 11996 5940 12000
rect 5876 11940 5880 11996
rect 5880 11940 5936 11996
rect 5936 11940 5940 11996
rect 5876 11936 5940 11940
rect 5956 11996 6020 12000
rect 5956 11940 5960 11996
rect 5960 11940 6016 11996
rect 6016 11940 6020 11996
rect 5956 11936 6020 11940
rect 6036 11996 6100 12000
rect 6036 11940 6040 11996
rect 6040 11940 6096 11996
rect 6096 11940 6100 11996
rect 6036 11936 6100 11940
rect 36516 11996 36580 12000
rect 36516 11940 36520 11996
rect 36520 11940 36576 11996
rect 36576 11940 36580 11996
rect 36516 11936 36580 11940
rect 36596 11996 36660 12000
rect 36596 11940 36600 11996
rect 36600 11940 36656 11996
rect 36656 11940 36660 11996
rect 36596 11936 36660 11940
rect 36676 11996 36740 12000
rect 36676 11940 36680 11996
rect 36680 11940 36736 11996
rect 36736 11940 36740 11996
rect 36676 11936 36740 11940
rect 36756 11996 36820 12000
rect 36756 11940 36760 11996
rect 36760 11940 36816 11996
rect 36816 11940 36820 11996
rect 36756 11936 36820 11940
rect 67236 11996 67300 12000
rect 67236 11940 67240 11996
rect 67240 11940 67296 11996
rect 67296 11940 67300 11996
rect 67236 11936 67300 11940
rect 67316 11996 67380 12000
rect 67316 11940 67320 11996
rect 67320 11940 67376 11996
rect 67376 11940 67380 11996
rect 67316 11936 67380 11940
rect 67396 11996 67460 12000
rect 67396 11940 67400 11996
rect 67400 11940 67456 11996
rect 67456 11940 67460 11996
rect 67396 11936 67460 11940
rect 67476 11996 67540 12000
rect 67476 11940 67480 11996
rect 67480 11940 67536 11996
rect 67536 11940 67540 11996
rect 67476 11936 67540 11940
rect 5136 11452 5200 11456
rect 5136 11396 5140 11452
rect 5140 11396 5196 11452
rect 5196 11396 5200 11452
rect 5136 11392 5200 11396
rect 5216 11452 5280 11456
rect 5216 11396 5220 11452
rect 5220 11396 5276 11452
rect 5276 11396 5280 11452
rect 5216 11392 5280 11396
rect 5296 11452 5360 11456
rect 5296 11396 5300 11452
rect 5300 11396 5356 11452
rect 5356 11396 5360 11452
rect 5296 11392 5360 11396
rect 5376 11452 5440 11456
rect 5376 11396 5380 11452
rect 5380 11396 5436 11452
rect 5436 11396 5440 11452
rect 5376 11392 5440 11396
rect 35856 11452 35920 11456
rect 35856 11396 35860 11452
rect 35860 11396 35916 11452
rect 35916 11396 35920 11452
rect 35856 11392 35920 11396
rect 35936 11452 36000 11456
rect 35936 11396 35940 11452
rect 35940 11396 35996 11452
rect 35996 11396 36000 11452
rect 35936 11392 36000 11396
rect 36016 11452 36080 11456
rect 36016 11396 36020 11452
rect 36020 11396 36076 11452
rect 36076 11396 36080 11452
rect 36016 11392 36080 11396
rect 36096 11452 36160 11456
rect 36096 11396 36100 11452
rect 36100 11396 36156 11452
rect 36156 11396 36160 11452
rect 36096 11392 36160 11396
rect 66576 11452 66640 11456
rect 66576 11396 66580 11452
rect 66580 11396 66636 11452
rect 66636 11396 66640 11452
rect 66576 11392 66640 11396
rect 66656 11452 66720 11456
rect 66656 11396 66660 11452
rect 66660 11396 66716 11452
rect 66716 11396 66720 11452
rect 66656 11392 66720 11396
rect 66736 11452 66800 11456
rect 66736 11396 66740 11452
rect 66740 11396 66796 11452
rect 66796 11396 66800 11452
rect 66736 11392 66800 11396
rect 66816 11452 66880 11456
rect 66816 11396 66820 11452
rect 66820 11396 66876 11452
rect 66876 11396 66880 11452
rect 66816 11392 66880 11396
rect 5796 10908 5860 10912
rect 5796 10852 5800 10908
rect 5800 10852 5856 10908
rect 5856 10852 5860 10908
rect 5796 10848 5860 10852
rect 5876 10908 5940 10912
rect 5876 10852 5880 10908
rect 5880 10852 5936 10908
rect 5936 10852 5940 10908
rect 5876 10848 5940 10852
rect 5956 10908 6020 10912
rect 5956 10852 5960 10908
rect 5960 10852 6016 10908
rect 6016 10852 6020 10908
rect 5956 10848 6020 10852
rect 6036 10908 6100 10912
rect 6036 10852 6040 10908
rect 6040 10852 6096 10908
rect 6096 10852 6100 10908
rect 6036 10848 6100 10852
rect 36516 10908 36580 10912
rect 36516 10852 36520 10908
rect 36520 10852 36576 10908
rect 36576 10852 36580 10908
rect 36516 10848 36580 10852
rect 36596 10908 36660 10912
rect 36596 10852 36600 10908
rect 36600 10852 36656 10908
rect 36656 10852 36660 10908
rect 36596 10848 36660 10852
rect 36676 10908 36740 10912
rect 36676 10852 36680 10908
rect 36680 10852 36736 10908
rect 36736 10852 36740 10908
rect 36676 10848 36740 10852
rect 36756 10908 36820 10912
rect 36756 10852 36760 10908
rect 36760 10852 36816 10908
rect 36816 10852 36820 10908
rect 36756 10848 36820 10852
rect 67236 10908 67300 10912
rect 67236 10852 67240 10908
rect 67240 10852 67296 10908
rect 67296 10852 67300 10908
rect 67236 10848 67300 10852
rect 67316 10908 67380 10912
rect 67316 10852 67320 10908
rect 67320 10852 67376 10908
rect 67376 10852 67380 10908
rect 67316 10848 67380 10852
rect 67396 10908 67460 10912
rect 67396 10852 67400 10908
rect 67400 10852 67456 10908
rect 67456 10852 67460 10908
rect 67396 10848 67460 10852
rect 67476 10908 67540 10912
rect 67476 10852 67480 10908
rect 67480 10852 67536 10908
rect 67536 10852 67540 10908
rect 67476 10848 67540 10852
rect 5136 10364 5200 10368
rect 5136 10308 5140 10364
rect 5140 10308 5196 10364
rect 5196 10308 5200 10364
rect 5136 10304 5200 10308
rect 5216 10364 5280 10368
rect 5216 10308 5220 10364
rect 5220 10308 5276 10364
rect 5276 10308 5280 10364
rect 5216 10304 5280 10308
rect 5296 10364 5360 10368
rect 5296 10308 5300 10364
rect 5300 10308 5356 10364
rect 5356 10308 5360 10364
rect 5296 10304 5360 10308
rect 5376 10364 5440 10368
rect 5376 10308 5380 10364
rect 5380 10308 5436 10364
rect 5436 10308 5440 10364
rect 5376 10304 5440 10308
rect 35856 10364 35920 10368
rect 35856 10308 35860 10364
rect 35860 10308 35916 10364
rect 35916 10308 35920 10364
rect 35856 10304 35920 10308
rect 35936 10364 36000 10368
rect 35936 10308 35940 10364
rect 35940 10308 35996 10364
rect 35996 10308 36000 10364
rect 35936 10304 36000 10308
rect 36016 10364 36080 10368
rect 36016 10308 36020 10364
rect 36020 10308 36076 10364
rect 36076 10308 36080 10364
rect 36016 10304 36080 10308
rect 36096 10364 36160 10368
rect 36096 10308 36100 10364
rect 36100 10308 36156 10364
rect 36156 10308 36160 10364
rect 36096 10304 36160 10308
rect 66576 10364 66640 10368
rect 66576 10308 66580 10364
rect 66580 10308 66636 10364
rect 66636 10308 66640 10364
rect 66576 10304 66640 10308
rect 66656 10364 66720 10368
rect 66656 10308 66660 10364
rect 66660 10308 66716 10364
rect 66716 10308 66720 10364
rect 66656 10304 66720 10308
rect 66736 10364 66800 10368
rect 66736 10308 66740 10364
rect 66740 10308 66796 10364
rect 66796 10308 66800 10364
rect 66736 10304 66800 10308
rect 66816 10364 66880 10368
rect 66816 10308 66820 10364
rect 66820 10308 66876 10364
rect 66876 10308 66880 10364
rect 66816 10304 66880 10308
rect 5796 9820 5860 9824
rect 5796 9764 5800 9820
rect 5800 9764 5856 9820
rect 5856 9764 5860 9820
rect 5796 9760 5860 9764
rect 5876 9820 5940 9824
rect 5876 9764 5880 9820
rect 5880 9764 5936 9820
rect 5936 9764 5940 9820
rect 5876 9760 5940 9764
rect 5956 9820 6020 9824
rect 5956 9764 5960 9820
rect 5960 9764 6016 9820
rect 6016 9764 6020 9820
rect 5956 9760 6020 9764
rect 6036 9820 6100 9824
rect 6036 9764 6040 9820
rect 6040 9764 6096 9820
rect 6096 9764 6100 9820
rect 6036 9760 6100 9764
rect 36516 9820 36580 9824
rect 36516 9764 36520 9820
rect 36520 9764 36576 9820
rect 36576 9764 36580 9820
rect 36516 9760 36580 9764
rect 36596 9820 36660 9824
rect 36596 9764 36600 9820
rect 36600 9764 36656 9820
rect 36656 9764 36660 9820
rect 36596 9760 36660 9764
rect 36676 9820 36740 9824
rect 36676 9764 36680 9820
rect 36680 9764 36736 9820
rect 36736 9764 36740 9820
rect 36676 9760 36740 9764
rect 36756 9820 36820 9824
rect 36756 9764 36760 9820
rect 36760 9764 36816 9820
rect 36816 9764 36820 9820
rect 36756 9760 36820 9764
rect 67236 9820 67300 9824
rect 67236 9764 67240 9820
rect 67240 9764 67296 9820
rect 67296 9764 67300 9820
rect 67236 9760 67300 9764
rect 67316 9820 67380 9824
rect 67316 9764 67320 9820
rect 67320 9764 67376 9820
rect 67376 9764 67380 9820
rect 67316 9760 67380 9764
rect 67396 9820 67460 9824
rect 67396 9764 67400 9820
rect 67400 9764 67456 9820
rect 67456 9764 67460 9820
rect 67396 9760 67460 9764
rect 67476 9820 67540 9824
rect 67476 9764 67480 9820
rect 67480 9764 67536 9820
rect 67536 9764 67540 9820
rect 67476 9760 67540 9764
rect 5136 9276 5200 9280
rect 5136 9220 5140 9276
rect 5140 9220 5196 9276
rect 5196 9220 5200 9276
rect 5136 9216 5200 9220
rect 5216 9276 5280 9280
rect 5216 9220 5220 9276
rect 5220 9220 5276 9276
rect 5276 9220 5280 9276
rect 5216 9216 5280 9220
rect 5296 9276 5360 9280
rect 5296 9220 5300 9276
rect 5300 9220 5356 9276
rect 5356 9220 5360 9276
rect 5296 9216 5360 9220
rect 5376 9276 5440 9280
rect 5376 9220 5380 9276
rect 5380 9220 5436 9276
rect 5436 9220 5440 9276
rect 5376 9216 5440 9220
rect 35856 9276 35920 9280
rect 35856 9220 35860 9276
rect 35860 9220 35916 9276
rect 35916 9220 35920 9276
rect 35856 9216 35920 9220
rect 35936 9276 36000 9280
rect 35936 9220 35940 9276
rect 35940 9220 35996 9276
rect 35996 9220 36000 9276
rect 35936 9216 36000 9220
rect 36016 9276 36080 9280
rect 36016 9220 36020 9276
rect 36020 9220 36076 9276
rect 36076 9220 36080 9276
rect 36016 9216 36080 9220
rect 36096 9276 36160 9280
rect 36096 9220 36100 9276
rect 36100 9220 36156 9276
rect 36156 9220 36160 9276
rect 36096 9216 36160 9220
rect 66576 9276 66640 9280
rect 66576 9220 66580 9276
rect 66580 9220 66636 9276
rect 66636 9220 66640 9276
rect 66576 9216 66640 9220
rect 66656 9276 66720 9280
rect 66656 9220 66660 9276
rect 66660 9220 66716 9276
rect 66716 9220 66720 9276
rect 66656 9216 66720 9220
rect 66736 9276 66800 9280
rect 66736 9220 66740 9276
rect 66740 9220 66796 9276
rect 66796 9220 66800 9276
rect 66736 9216 66800 9220
rect 66816 9276 66880 9280
rect 66816 9220 66820 9276
rect 66820 9220 66876 9276
rect 66876 9220 66880 9276
rect 66816 9216 66880 9220
rect 5796 8732 5860 8736
rect 5796 8676 5800 8732
rect 5800 8676 5856 8732
rect 5856 8676 5860 8732
rect 5796 8672 5860 8676
rect 5876 8732 5940 8736
rect 5876 8676 5880 8732
rect 5880 8676 5936 8732
rect 5936 8676 5940 8732
rect 5876 8672 5940 8676
rect 5956 8732 6020 8736
rect 5956 8676 5960 8732
rect 5960 8676 6016 8732
rect 6016 8676 6020 8732
rect 5956 8672 6020 8676
rect 6036 8732 6100 8736
rect 6036 8676 6040 8732
rect 6040 8676 6096 8732
rect 6096 8676 6100 8732
rect 6036 8672 6100 8676
rect 36516 8732 36580 8736
rect 36516 8676 36520 8732
rect 36520 8676 36576 8732
rect 36576 8676 36580 8732
rect 36516 8672 36580 8676
rect 36596 8732 36660 8736
rect 36596 8676 36600 8732
rect 36600 8676 36656 8732
rect 36656 8676 36660 8732
rect 36596 8672 36660 8676
rect 36676 8732 36740 8736
rect 36676 8676 36680 8732
rect 36680 8676 36736 8732
rect 36736 8676 36740 8732
rect 36676 8672 36740 8676
rect 36756 8732 36820 8736
rect 36756 8676 36760 8732
rect 36760 8676 36816 8732
rect 36816 8676 36820 8732
rect 36756 8672 36820 8676
rect 67236 8732 67300 8736
rect 67236 8676 67240 8732
rect 67240 8676 67296 8732
rect 67296 8676 67300 8732
rect 67236 8672 67300 8676
rect 67316 8732 67380 8736
rect 67316 8676 67320 8732
rect 67320 8676 67376 8732
rect 67376 8676 67380 8732
rect 67316 8672 67380 8676
rect 67396 8732 67460 8736
rect 67396 8676 67400 8732
rect 67400 8676 67456 8732
rect 67456 8676 67460 8732
rect 67396 8672 67460 8676
rect 67476 8732 67540 8736
rect 67476 8676 67480 8732
rect 67480 8676 67536 8732
rect 67536 8676 67540 8732
rect 67476 8672 67540 8676
rect 5136 8188 5200 8192
rect 5136 8132 5140 8188
rect 5140 8132 5196 8188
rect 5196 8132 5200 8188
rect 5136 8128 5200 8132
rect 5216 8188 5280 8192
rect 5216 8132 5220 8188
rect 5220 8132 5276 8188
rect 5276 8132 5280 8188
rect 5216 8128 5280 8132
rect 5296 8188 5360 8192
rect 5296 8132 5300 8188
rect 5300 8132 5356 8188
rect 5356 8132 5360 8188
rect 5296 8128 5360 8132
rect 5376 8188 5440 8192
rect 5376 8132 5380 8188
rect 5380 8132 5436 8188
rect 5436 8132 5440 8188
rect 5376 8128 5440 8132
rect 35856 8188 35920 8192
rect 35856 8132 35860 8188
rect 35860 8132 35916 8188
rect 35916 8132 35920 8188
rect 35856 8128 35920 8132
rect 35936 8188 36000 8192
rect 35936 8132 35940 8188
rect 35940 8132 35996 8188
rect 35996 8132 36000 8188
rect 35936 8128 36000 8132
rect 36016 8188 36080 8192
rect 36016 8132 36020 8188
rect 36020 8132 36076 8188
rect 36076 8132 36080 8188
rect 36016 8128 36080 8132
rect 36096 8188 36160 8192
rect 36096 8132 36100 8188
rect 36100 8132 36156 8188
rect 36156 8132 36160 8188
rect 36096 8128 36160 8132
rect 66576 8188 66640 8192
rect 66576 8132 66580 8188
rect 66580 8132 66636 8188
rect 66636 8132 66640 8188
rect 66576 8128 66640 8132
rect 66656 8188 66720 8192
rect 66656 8132 66660 8188
rect 66660 8132 66716 8188
rect 66716 8132 66720 8188
rect 66656 8128 66720 8132
rect 66736 8188 66800 8192
rect 66736 8132 66740 8188
rect 66740 8132 66796 8188
rect 66796 8132 66800 8188
rect 66736 8128 66800 8132
rect 66816 8188 66880 8192
rect 66816 8132 66820 8188
rect 66820 8132 66876 8188
rect 66876 8132 66880 8188
rect 66816 8128 66880 8132
rect 5796 7644 5860 7648
rect 5796 7588 5800 7644
rect 5800 7588 5856 7644
rect 5856 7588 5860 7644
rect 5796 7584 5860 7588
rect 5876 7644 5940 7648
rect 5876 7588 5880 7644
rect 5880 7588 5936 7644
rect 5936 7588 5940 7644
rect 5876 7584 5940 7588
rect 5956 7644 6020 7648
rect 5956 7588 5960 7644
rect 5960 7588 6016 7644
rect 6016 7588 6020 7644
rect 5956 7584 6020 7588
rect 6036 7644 6100 7648
rect 6036 7588 6040 7644
rect 6040 7588 6096 7644
rect 6096 7588 6100 7644
rect 6036 7584 6100 7588
rect 36516 7644 36580 7648
rect 36516 7588 36520 7644
rect 36520 7588 36576 7644
rect 36576 7588 36580 7644
rect 36516 7584 36580 7588
rect 36596 7644 36660 7648
rect 36596 7588 36600 7644
rect 36600 7588 36656 7644
rect 36656 7588 36660 7644
rect 36596 7584 36660 7588
rect 36676 7644 36740 7648
rect 36676 7588 36680 7644
rect 36680 7588 36736 7644
rect 36736 7588 36740 7644
rect 36676 7584 36740 7588
rect 36756 7644 36820 7648
rect 36756 7588 36760 7644
rect 36760 7588 36816 7644
rect 36816 7588 36820 7644
rect 36756 7584 36820 7588
rect 67236 7644 67300 7648
rect 67236 7588 67240 7644
rect 67240 7588 67296 7644
rect 67296 7588 67300 7644
rect 67236 7584 67300 7588
rect 67316 7644 67380 7648
rect 67316 7588 67320 7644
rect 67320 7588 67376 7644
rect 67376 7588 67380 7644
rect 67316 7584 67380 7588
rect 67396 7644 67460 7648
rect 67396 7588 67400 7644
rect 67400 7588 67456 7644
rect 67456 7588 67460 7644
rect 67396 7584 67460 7588
rect 67476 7644 67540 7648
rect 67476 7588 67480 7644
rect 67480 7588 67536 7644
rect 67536 7588 67540 7644
rect 67476 7584 67540 7588
rect 5136 7100 5200 7104
rect 5136 7044 5140 7100
rect 5140 7044 5196 7100
rect 5196 7044 5200 7100
rect 5136 7040 5200 7044
rect 5216 7100 5280 7104
rect 5216 7044 5220 7100
rect 5220 7044 5276 7100
rect 5276 7044 5280 7100
rect 5216 7040 5280 7044
rect 5296 7100 5360 7104
rect 5296 7044 5300 7100
rect 5300 7044 5356 7100
rect 5356 7044 5360 7100
rect 5296 7040 5360 7044
rect 5376 7100 5440 7104
rect 5376 7044 5380 7100
rect 5380 7044 5436 7100
rect 5436 7044 5440 7100
rect 5376 7040 5440 7044
rect 35856 7100 35920 7104
rect 35856 7044 35860 7100
rect 35860 7044 35916 7100
rect 35916 7044 35920 7100
rect 35856 7040 35920 7044
rect 35936 7100 36000 7104
rect 35936 7044 35940 7100
rect 35940 7044 35996 7100
rect 35996 7044 36000 7100
rect 35936 7040 36000 7044
rect 36016 7100 36080 7104
rect 36016 7044 36020 7100
rect 36020 7044 36076 7100
rect 36076 7044 36080 7100
rect 36016 7040 36080 7044
rect 36096 7100 36160 7104
rect 36096 7044 36100 7100
rect 36100 7044 36156 7100
rect 36156 7044 36160 7100
rect 36096 7040 36160 7044
rect 66576 7100 66640 7104
rect 66576 7044 66580 7100
rect 66580 7044 66636 7100
rect 66636 7044 66640 7100
rect 66576 7040 66640 7044
rect 66656 7100 66720 7104
rect 66656 7044 66660 7100
rect 66660 7044 66716 7100
rect 66716 7044 66720 7100
rect 66656 7040 66720 7044
rect 66736 7100 66800 7104
rect 66736 7044 66740 7100
rect 66740 7044 66796 7100
rect 66796 7044 66800 7100
rect 66736 7040 66800 7044
rect 66816 7100 66880 7104
rect 66816 7044 66820 7100
rect 66820 7044 66876 7100
rect 66876 7044 66880 7100
rect 66816 7040 66880 7044
rect 5796 6556 5860 6560
rect 5796 6500 5800 6556
rect 5800 6500 5856 6556
rect 5856 6500 5860 6556
rect 5796 6496 5860 6500
rect 5876 6556 5940 6560
rect 5876 6500 5880 6556
rect 5880 6500 5936 6556
rect 5936 6500 5940 6556
rect 5876 6496 5940 6500
rect 5956 6556 6020 6560
rect 5956 6500 5960 6556
rect 5960 6500 6016 6556
rect 6016 6500 6020 6556
rect 5956 6496 6020 6500
rect 6036 6556 6100 6560
rect 6036 6500 6040 6556
rect 6040 6500 6096 6556
rect 6096 6500 6100 6556
rect 6036 6496 6100 6500
rect 36516 6556 36580 6560
rect 36516 6500 36520 6556
rect 36520 6500 36576 6556
rect 36576 6500 36580 6556
rect 36516 6496 36580 6500
rect 36596 6556 36660 6560
rect 36596 6500 36600 6556
rect 36600 6500 36656 6556
rect 36656 6500 36660 6556
rect 36596 6496 36660 6500
rect 36676 6556 36740 6560
rect 36676 6500 36680 6556
rect 36680 6500 36736 6556
rect 36736 6500 36740 6556
rect 36676 6496 36740 6500
rect 36756 6556 36820 6560
rect 36756 6500 36760 6556
rect 36760 6500 36816 6556
rect 36816 6500 36820 6556
rect 36756 6496 36820 6500
rect 67236 6556 67300 6560
rect 67236 6500 67240 6556
rect 67240 6500 67296 6556
rect 67296 6500 67300 6556
rect 67236 6496 67300 6500
rect 67316 6556 67380 6560
rect 67316 6500 67320 6556
rect 67320 6500 67376 6556
rect 67376 6500 67380 6556
rect 67316 6496 67380 6500
rect 67396 6556 67460 6560
rect 67396 6500 67400 6556
rect 67400 6500 67456 6556
rect 67456 6500 67460 6556
rect 67396 6496 67460 6500
rect 67476 6556 67540 6560
rect 67476 6500 67480 6556
rect 67480 6500 67536 6556
rect 67536 6500 67540 6556
rect 67476 6496 67540 6500
rect 5136 6012 5200 6016
rect 5136 5956 5140 6012
rect 5140 5956 5196 6012
rect 5196 5956 5200 6012
rect 5136 5952 5200 5956
rect 5216 6012 5280 6016
rect 5216 5956 5220 6012
rect 5220 5956 5276 6012
rect 5276 5956 5280 6012
rect 5216 5952 5280 5956
rect 5296 6012 5360 6016
rect 5296 5956 5300 6012
rect 5300 5956 5356 6012
rect 5356 5956 5360 6012
rect 5296 5952 5360 5956
rect 5376 6012 5440 6016
rect 5376 5956 5380 6012
rect 5380 5956 5436 6012
rect 5436 5956 5440 6012
rect 5376 5952 5440 5956
rect 35856 6012 35920 6016
rect 35856 5956 35860 6012
rect 35860 5956 35916 6012
rect 35916 5956 35920 6012
rect 35856 5952 35920 5956
rect 35936 6012 36000 6016
rect 35936 5956 35940 6012
rect 35940 5956 35996 6012
rect 35996 5956 36000 6012
rect 35936 5952 36000 5956
rect 36016 6012 36080 6016
rect 36016 5956 36020 6012
rect 36020 5956 36076 6012
rect 36076 5956 36080 6012
rect 36016 5952 36080 5956
rect 36096 6012 36160 6016
rect 36096 5956 36100 6012
rect 36100 5956 36156 6012
rect 36156 5956 36160 6012
rect 36096 5952 36160 5956
rect 66576 6012 66640 6016
rect 66576 5956 66580 6012
rect 66580 5956 66636 6012
rect 66636 5956 66640 6012
rect 66576 5952 66640 5956
rect 66656 6012 66720 6016
rect 66656 5956 66660 6012
rect 66660 5956 66716 6012
rect 66716 5956 66720 6012
rect 66656 5952 66720 5956
rect 66736 6012 66800 6016
rect 66736 5956 66740 6012
rect 66740 5956 66796 6012
rect 66796 5956 66800 6012
rect 66736 5952 66800 5956
rect 66816 6012 66880 6016
rect 66816 5956 66820 6012
rect 66820 5956 66876 6012
rect 66876 5956 66880 6012
rect 66816 5952 66880 5956
rect 5796 5468 5860 5472
rect 5796 5412 5800 5468
rect 5800 5412 5856 5468
rect 5856 5412 5860 5468
rect 5796 5408 5860 5412
rect 5876 5468 5940 5472
rect 5876 5412 5880 5468
rect 5880 5412 5936 5468
rect 5936 5412 5940 5468
rect 5876 5408 5940 5412
rect 5956 5468 6020 5472
rect 5956 5412 5960 5468
rect 5960 5412 6016 5468
rect 6016 5412 6020 5468
rect 5956 5408 6020 5412
rect 6036 5468 6100 5472
rect 6036 5412 6040 5468
rect 6040 5412 6096 5468
rect 6096 5412 6100 5468
rect 6036 5408 6100 5412
rect 36516 5468 36580 5472
rect 36516 5412 36520 5468
rect 36520 5412 36576 5468
rect 36576 5412 36580 5468
rect 36516 5408 36580 5412
rect 36596 5468 36660 5472
rect 36596 5412 36600 5468
rect 36600 5412 36656 5468
rect 36656 5412 36660 5468
rect 36596 5408 36660 5412
rect 36676 5468 36740 5472
rect 36676 5412 36680 5468
rect 36680 5412 36736 5468
rect 36736 5412 36740 5468
rect 36676 5408 36740 5412
rect 36756 5468 36820 5472
rect 36756 5412 36760 5468
rect 36760 5412 36816 5468
rect 36816 5412 36820 5468
rect 36756 5408 36820 5412
rect 67236 5468 67300 5472
rect 67236 5412 67240 5468
rect 67240 5412 67296 5468
rect 67296 5412 67300 5468
rect 67236 5408 67300 5412
rect 67316 5468 67380 5472
rect 67316 5412 67320 5468
rect 67320 5412 67376 5468
rect 67376 5412 67380 5468
rect 67316 5408 67380 5412
rect 67396 5468 67460 5472
rect 67396 5412 67400 5468
rect 67400 5412 67456 5468
rect 67456 5412 67460 5468
rect 67396 5408 67460 5412
rect 67476 5468 67540 5472
rect 67476 5412 67480 5468
rect 67480 5412 67536 5468
rect 67536 5412 67540 5468
rect 67476 5408 67540 5412
rect 5136 4924 5200 4928
rect 5136 4868 5140 4924
rect 5140 4868 5196 4924
rect 5196 4868 5200 4924
rect 5136 4864 5200 4868
rect 5216 4924 5280 4928
rect 5216 4868 5220 4924
rect 5220 4868 5276 4924
rect 5276 4868 5280 4924
rect 5216 4864 5280 4868
rect 5296 4924 5360 4928
rect 5296 4868 5300 4924
rect 5300 4868 5356 4924
rect 5356 4868 5360 4924
rect 5296 4864 5360 4868
rect 5376 4924 5440 4928
rect 5376 4868 5380 4924
rect 5380 4868 5436 4924
rect 5436 4868 5440 4924
rect 5376 4864 5440 4868
rect 35856 4924 35920 4928
rect 35856 4868 35860 4924
rect 35860 4868 35916 4924
rect 35916 4868 35920 4924
rect 35856 4864 35920 4868
rect 35936 4924 36000 4928
rect 35936 4868 35940 4924
rect 35940 4868 35996 4924
rect 35996 4868 36000 4924
rect 35936 4864 36000 4868
rect 36016 4924 36080 4928
rect 36016 4868 36020 4924
rect 36020 4868 36076 4924
rect 36076 4868 36080 4924
rect 36016 4864 36080 4868
rect 36096 4924 36160 4928
rect 36096 4868 36100 4924
rect 36100 4868 36156 4924
rect 36156 4868 36160 4924
rect 36096 4864 36160 4868
rect 66576 4924 66640 4928
rect 66576 4868 66580 4924
rect 66580 4868 66636 4924
rect 66636 4868 66640 4924
rect 66576 4864 66640 4868
rect 66656 4924 66720 4928
rect 66656 4868 66660 4924
rect 66660 4868 66716 4924
rect 66716 4868 66720 4924
rect 66656 4864 66720 4868
rect 66736 4924 66800 4928
rect 66736 4868 66740 4924
rect 66740 4868 66796 4924
rect 66796 4868 66800 4924
rect 66736 4864 66800 4868
rect 66816 4924 66880 4928
rect 66816 4868 66820 4924
rect 66820 4868 66876 4924
rect 66876 4868 66880 4924
rect 66816 4864 66880 4868
rect 5796 4380 5860 4384
rect 5796 4324 5800 4380
rect 5800 4324 5856 4380
rect 5856 4324 5860 4380
rect 5796 4320 5860 4324
rect 5876 4380 5940 4384
rect 5876 4324 5880 4380
rect 5880 4324 5936 4380
rect 5936 4324 5940 4380
rect 5876 4320 5940 4324
rect 5956 4380 6020 4384
rect 5956 4324 5960 4380
rect 5960 4324 6016 4380
rect 6016 4324 6020 4380
rect 5956 4320 6020 4324
rect 6036 4380 6100 4384
rect 6036 4324 6040 4380
rect 6040 4324 6096 4380
rect 6096 4324 6100 4380
rect 6036 4320 6100 4324
rect 36516 4380 36580 4384
rect 36516 4324 36520 4380
rect 36520 4324 36576 4380
rect 36576 4324 36580 4380
rect 36516 4320 36580 4324
rect 36596 4380 36660 4384
rect 36596 4324 36600 4380
rect 36600 4324 36656 4380
rect 36656 4324 36660 4380
rect 36596 4320 36660 4324
rect 36676 4380 36740 4384
rect 36676 4324 36680 4380
rect 36680 4324 36736 4380
rect 36736 4324 36740 4380
rect 36676 4320 36740 4324
rect 36756 4380 36820 4384
rect 36756 4324 36760 4380
rect 36760 4324 36816 4380
rect 36816 4324 36820 4380
rect 36756 4320 36820 4324
rect 67236 4380 67300 4384
rect 67236 4324 67240 4380
rect 67240 4324 67296 4380
rect 67296 4324 67300 4380
rect 67236 4320 67300 4324
rect 67316 4380 67380 4384
rect 67316 4324 67320 4380
rect 67320 4324 67376 4380
rect 67376 4324 67380 4380
rect 67316 4320 67380 4324
rect 67396 4380 67460 4384
rect 67396 4324 67400 4380
rect 67400 4324 67456 4380
rect 67456 4324 67460 4380
rect 67396 4320 67460 4324
rect 67476 4380 67540 4384
rect 67476 4324 67480 4380
rect 67480 4324 67536 4380
rect 67536 4324 67540 4380
rect 67476 4320 67540 4324
rect 5136 3836 5200 3840
rect 5136 3780 5140 3836
rect 5140 3780 5196 3836
rect 5196 3780 5200 3836
rect 5136 3776 5200 3780
rect 5216 3836 5280 3840
rect 5216 3780 5220 3836
rect 5220 3780 5276 3836
rect 5276 3780 5280 3836
rect 5216 3776 5280 3780
rect 5296 3836 5360 3840
rect 5296 3780 5300 3836
rect 5300 3780 5356 3836
rect 5356 3780 5360 3836
rect 5296 3776 5360 3780
rect 5376 3836 5440 3840
rect 5376 3780 5380 3836
rect 5380 3780 5436 3836
rect 5436 3780 5440 3836
rect 5376 3776 5440 3780
rect 35856 3836 35920 3840
rect 35856 3780 35860 3836
rect 35860 3780 35916 3836
rect 35916 3780 35920 3836
rect 35856 3776 35920 3780
rect 35936 3836 36000 3840
rect 35936 3780 35940 3836
rect 35940 3780 35996 3836
rect 35996 3780 36000 3836
rect 35936 3776 36000 3780
rect 36016 3836 36080 3840
rect 36016 3780 36020 3836
rect 36020 3780 36076 3836
rect 36076 3780 36080 3836
rect 36016 3776 36080 3780
rect 36096 3836 36160 3840
rect 36096 3780 36100 3836
rect 36100 3780 36156 3836
rect 36156 3780 36160 3836
rect 36096 3776 36160 3780
rect 66576 3836 66640 3840
rect 66576 3780 66580 3836
rect 66580 3780 66636 3836
rect 66636 3780 66640 3836
rect 66576 3776 66640 3780
rect 66656 3836 66720 3840
rect 66656 3780 66660 3836
rect 66660 3780 66716 3836
rect 66716 3780 66720 3836
rect 66656 3776 66720 3780
rect 66736 3836 66800 3840
rect 66736 3780 66740 3836
rect 66740 3780 66796 3836
rect 66796 3780 66800 3836
rect 66736 3776 66800 3780
rect 66816 3836 66880 3840
rect 66816 3780 66820 3836
rect 66820 3780 66876 3836
rect 66876 3780 66880 3836
rect 66816 3776 66880 3780
rect 5796 3292 5860 3296
rect 5796 3236 5800 3292
rect 5800 3236 5856 3292
rect 5856 3236 5860 3292
rect 5796 3232 5860 3236
rect 5876 3292 5940 3296
rect 5876 3236 5880 3292
rect 5880 3236 5936 3292
rect 5936 3236 5940 3292
rect 5876 3232 5940 3236
rect 5956 3292 6020 3296
rect 5956 3236 5960 3292
rect 5960 3236 6016 3292
rect 6016 3236 6020 3292
rect 5956 3232 6020 3236
rect 6036 3292 6100 3296
rect 6036 3236 6040 3292
rect 6040 3236 6096 3292
rect 6096 3236 6100 3292
rect 6036 3232 6100 3236
rect 36516 3292 36580 3296
rect 36516 3236 36520 3292
rect 36520 3236 36576 3292
rect 36576 3236 36580 3292
rect 36516 3232 36580 3236
rect 36596 3292 36660 3296
rect 36596 3236 36600 3292
rect 36600 3236 36656 3292
rect 36656 3236 36660 3292
rect 36596 3232 36660 3236
rect 36676 3292 36740 3296
rect 36676 3236 36680 3292
rect 36680 3236 36736 3292
rect 36736 3236 36740 3292
rect 36676 3232 36740 3236
rect 36756 3292 36820 3296
rect 36756 3236 36760 3292
rect 36760 3236 36816 3292
rect 36816 3236 36820 3292
rect 36756 3232 36820 3236
rect 67236 3292 67300 3296
rect 67236 3236 67240 3292
rect 67240 3236 67296 3292
rect 67296 3236 67300 3292
rect 67236 3232 67300 3236
rect 67316 3292 67380 3296
rect 67316 3236 67320 3292
rect 67320 3236 67376 3292
rect 67376 3236 67380 3292
rect 67316 3232 67380 3236
rect 67396 3292 67460 3296
rect 67396 3236 67400 3292
rect 67400 3236 67456 3292
rect 67456 3236 67460 3292
rect 67396 3232 67460 3236
rect 67476 3292 67540 3296
rect 67476 3236 67480 3292
rect 67480 3236 67536 3292
rect 67536 3236 67540 3292
rect 67476 3232 67540 3236
rect 5136 2748 5200 2752
rect 5136 2692 5140 2748
rect 5140 2692 5196 2748
rect 5196 2692 5200 2748
rect 5136 2688 5200 2692
rect 5216 2748 5280 2752
rect 5216 2692 5220 2748
rect 5220 2692 5276 2748
rect 5276 2692 5280 2748
rect 5216 2688 5280 2692
rect 5296 2748 5360 2752
rect 5296 2692 5300 2748
rect 5300 2692 5356 2748
rect 5356 2692 5360 2748
rect 5296 2688 5360 2692
rect 5376 2748 5440 2752
rect 5376 2692 5380 2748
rect 5380 2692 5436 2748
rect 5436 2692 5440 2748
rect 5376 2688 5440 2692
rect 35856 2748 35920 2752
rect 35856 2692 35860 2748
rect 35860 2692 35916 2748
rect 35916 2692 35920 2748
rect 35856 2688 35920 2692
rect 35936 2748 36000 2752
rect 35936 2692 35940 2748
rect 35940 2692 35996 2748
rect 35996 2692 36000 2748
rect 35936 2688 36000 2692
rect 36016 2748 36080 2752
rect 36016 2692 36020 2748
rect 36020 2692 36076 2748
rect 36076 2692 36080 2748
rect 36016 2688 36080 2692
rect 36096 2748 36160 2752
rect 36096 2692 36100 2748
rect 36100 2692 36156 2748
rect 36156 2692 36160 2748
rect 36096 2688 36160 2692
rect 66576 2748 66640 2752
rect 66576 2692 66580 2748
rect 66580 2692 66636 2748
rect 66636 2692 66640 2748
rect 66576 2688 66640 2692
rect 66656 2748 66720 2752
rect 66656 2692 66660 2748
rect 66660 2692 66716 2748
rect 66716 2692 66720 2748
rect 66656 2688 66720 2692
rect 66736 2748 66800 2752
rect 66736 2692 66740 2748
rect 66740 2692 66796 2748
rect 66796 2692 66800 2748
rect 66736 2688 66800 2692
rect 66816 2748 66880 2752
rect 66816 2692 66820 2748
rect 66820 2692 66876 2748
rect 66876 2692 66880 2748
rect 66816 2688 66880 2692
rect 5796 2204 5860 2208
rect 5796 2148 5800 2204
rect 5800 2148 5856 2204
rect 5856 2148 5860 2204
rect 5796 2144 5860 2148
rect 5876 2204 5940 2208
rect 5876 2148 5880 2204
rect 5880 2148 5936 2204
rect 5936 2148 5940 2204
rect 5876 2144 5940 2148
rect 5956 2204 6020 2208
rect 5956 2148 5960 2204
rect 5960 2148 6016 2204
rect 6016 2148 6020 2204
rect 5956 2144 6020 2148
rect 6036 2204 6100 2208
rect 6036 2148 6040 2204
rect 6040 2148 6096 2204
rect 6096 2148 6100 2204
rect 6036 2144 6100 2148
rect 36516 2204 36580 2208
rect 36516 2148 36520 2204
rect 36520 2148 36576 2204
rect 36576 2148 36580 2204
rect 36516 2144 36580 2148
rect 36596 2204 36660 2208
rect 36596 2148 36600 2204
rect 36600 2148 36656 2204
rect 36656 2148 36660 2204
rect 36596 2144 36660 2148
rect 36676 2204 36740 2208
rect 36676 2148 36680 2204
rect 36680 2148 36736 2204
rect 36736 2148 36740 2204
rect 36676 2144 36740 2148
rect 36756 2204 36820 2208
rect 36756 2148 36760 2204
rect 36760 2148 36816 2204
rect 36816 2148 36820 2204
rect 36756 2144 36820 2148
rect 67236 2204 67300 2208
rect 67236 2148 67240 2204
rect 67240 2148 67296 2204
rect 67296 2148 67300 2204
rect 67236 2144 67300 2148
rect 67316 2204 67380 2208
rect 67316 2148 67320 2204
rect 67320 2148 67376 2204
rect 67376 2148 67380 2204
rect 67316 2144 67380 2148
rect 67396 2204 67460 2208
rect 67396 2148 67400 2204
rect 67400 2148 67456 2204
rect 67456 2148 67460 2204
rect 67396 2144 67460 2148
rect 67476 2204 67540 2208
rect 67476 2148 67480 2204
rect 67480 2148 67536 2204
rect 67536 2148 67540 2204
rect 67476 2144 67540 2148
<< metal4 >>
rect 5128 77824 5448 77840
rect 5128 77760 5136 77824
rect 5200 77760 5216 77824
rect 5280 77760 5296 77824
rect 5360 77760 5376 77824
rect 5440 77760 5448 77824
rect 5128 76736 5448 77760
rect 5128 76672 5136 76736
rect 5200 76672 5216 76736
rect 5280 76672 5296 76736
rect 5360 76672 5376 76736
rect 5440 76672 5448 76736
rect 5128 75648 5448 76672
rect 5128 75584 5136 75648
rect 5200 75584 5216 75648
rect 5280 75584 5296 75648
rect 5360 75584 5376 75648
rect 5440 75584 5448 75648
rect 5128 74560 5448 75584
rect 5128 74496 5136 74560
rect 5200 74496 5216 74560
rect 5280 74496 5296 74560
rect 5360 74496 5376 74560
rect 5440 74496 5448 74560
rect 5128 73472 5448 74496
rect 5128 73408 5136 73472
rect 5200 73408 5216 73472
rect 5280 73408 5296 73472
rect 5360 73408 5376 73472
rect 5440 73408 5448 73472
rect 5128 72384 5448 73408
rect 5128 72320 5136 72384
rect 5200 72320 5216 72384
rect 5280 72320 5296 72384
rect 5360 72320 5376 72384
rect 5440 72320 5448 72384
rect 5128 71296 5448 72320
rect 5128 71232 5136 71296
rect 5200 71232 5216 71296
rect 5280 71232 5296 71296
rect 5360 71232 5376 71296
rect 5440 71232 5448 71296
rect 5128 70208 5448 71232
rect 5128 70144 5136 70208
rect 5200 70144 5216 70208
rect 5280 70144 5296 70208
rect 5360 70144 5376 70208
rect 5440 70144 5448 70208
rect 5128 69120 5448 70144
rect 5128 69056 5136 69120
rect 5200 69056 5216 69120
rect 5280 69056 5296 69120
rect 5360 69056 5376 69120
rect 5440 69056 5448 69120
rect 5128 68032 5448 69056
rect 5128 67968 5136 68032
rect 5200 67968 5216 68032
rect 5280 67968 5296 68032
rect 5360 67968 5376 68032
rect 5440 67968 5448 68032
rect 5128 66944 5448 67968
rect 5128 66880 5136 66944
rect 5200 66896 5216 66944
rect 5280 66896 5296 66944
rect 5360 66896 5376 66944
rect 5440 66880 5448 66944
rect 5128 66660 5170 66880
rect 5406 66660 5448 66880
rect 5128 65856 5448 66660
rect 5128 65792 5136 65856
rect 5200 65792 5216 65856
rect 5280 65792 5296 65856
rect 5360 65792 5376 65856
rect 5440 65792 5448 65856
rect 5128 64768 5448 65792
rect 5128 64704 5136 64768
rect 5200 64704 5216 64768
rect 5280 64704 5296 64768
rect 5360 64704 5376 64768
rect 5440 64704 5448 64768
rect 5128 63680 5448 64704
rect 5128 63616 5136 63680
rect 5200 63616 5216 63680
rect 5280 63616 5296 63680
rect 5360 63616 5376 63680
rect 5440 63616 5448 63680
rect 5128 62592 5448 63616
rect 5128 62528 5136 62592
rect 5200 62528 5216 62592
rect 5280 62528 5296 62592
rect 5360 62528 5376 62592
rect 5440 62528 5448 62592
rect 5128 61504 5448 62528
rect 5128 61440 5136 61504
rect 5200 61440 5216 61504
rect 5280 61440 5296 61504
rect 5360 61440 5376 61504
rect 5440 61440 5448 61504
rect 5128 60416 5448 61440
rect 5128 60352 5136 60416
rect 5200 60352 5216 60416
rect 5280 60352 5296 60416
rect 5360 60352 5376 60416
rect 5440 60352 5448 60416
rect 5128 59328 5448 60352
rect 5128 59264 5136 59328
rect 5200 59264 5216 59328
rect 5280 59264 5296 59328
rect 5360 59264 5376 59328
rect 5440 59264 5448 59328
rect 5128 58240 5448 59264
rect 5128 58176 5136 58240
rect 5200 58176 5216 58240
rect 5280 58176 5296 58240
rect 5360 58176 5376 58240
rect 5440 58176 5448 58240
rect 5128 57152 5448 58176
rect 5128 57088 5136 57152
rect 5200 57088 5216 57152
rect 5280 57088 5296 57152
rect 5360 57088 5376 57152
rect 5440 57088 5448 57152
rect 5128 56064 5448 57088
rect 5128 56000 5136 56064
rect 5200 56000 5216 56064
rect 5280 56000 5296 56064
rect 5360 56000 5376 56064
rect 5440 56000 5448 56064
rect 5128 54976 5448 56000
rect 5128 54912 5136 54976
rect 5200 54912 5216 54976
rect 5280 54912 5296 54976
rect 5360 54912 5376 54976
rect 5440 54912 5448 54976
rect 5128 53888 5448 54912
rect 5128 53824 5136 53888
rect 5200 53824 5216 53888
rect 5280 53824 5296 53888
rect 5360 53824 5376 53888
rect 5440 53824 5448 53888
rect 5128 52800 5448 53824
rect 5128 52736 5136 52800
rect 5200 52736 5216 52800
rect 5280 52736 5296 52800
rect 5360 52736 5376 52800
rect 5440 52736 5448 52800
rect 5128 51712 5448 52736
rect 5128 51648 5136 51712
rect 5200 51648 5216 51712
rect 5280 51648 5296 51712
rect 5360 51648 5376 51712
rect 5440 51648 5448 51712
rect 5128 50624 5448 51648
rect 5128 50560 5136 50624
rect 5200 50560 5216 50624
rect 5280 50560 5296 50624
rect 5360 50560 5376 50624
rect 5440 50560 5448 50624
rect 5128 49536 5448 50560
rect 5128 49472 5136 49536
rect 5200 49472 5216 49536
rect 5280 49472 5296 49536
rect 5360 49472 5376 49536
rect 5440 49472 5448 49536
rect 5128 48448 5448 49472
rect 5128 48384 5136 48448
rect 5200 48384 5216 48448
rect 5280 48384 5296 48448
rect 5360 48384 5376 48448
rect 5440 48384 5448 48448
rect 5128 47360 5448 48384
rect 5128 47296 5136 47360
rect 5200 47296 5216 47360
rect 5280 47296 5296 47360
rect 5360 47296 5376 47360
rect 5440 47296 5448 47360
rect 5128 46272 5448 47296
rect 5128 46208 5136 46272
rect 5200 46208 5216 46272
rect 5280 46208 5296 46272
rect 5360 46208 5376 46272
rect 5440 46208 5448 46272
rect 5128 45184 5448 46208
rect 5128 45120 5136 45184
rect 5200 45120 5216 45184
rect 5280 45120 5296 45184
rect 5360 45120 5376 45184
rect 5440 45120 5448 45184
rect 5128 44096 5448 45120
rect 5128 44032 5136 44096
rect 5200 44032 5216 44096
rect 5280 44032 5296 44096
rect 5360 44032 5376 44096
rect 5440 44032 5448 44096
rect 5128 43008 5448 44032
rect 5128 42944 5136 43008
rect 5200 42944 5216 43008
rect 5280 42944 5296 43008
rect 5360 42944 5376 43008
rect 5440 42944 5448 43008
rect 5128 41920 5448 42944
rect 5128 41856 5136 41920
rect 5200 41856 5216 41920
rect 5280 41856 5296 41920
rect 5360 41856 5376 41920
rect 5440 41856 5448 41920
rect 5128 40832 5448 41856
rect 5128 40768 5136 40832
rect 5200 40768 5216 40832
rect 5280 40768 5296 40832
rect 5360 40768 5376 40832
rect 5440 40768 5448 40832
rect 5128 39744 5448 40768
rect 5128 39680 5136 39744
rect 5200 39680 5216 39744
rect 5280 39680 5296 39744
rect 5360 39680 5376 39744
rect 5440 39680 5448 39744
rect 5128 38656 5448 39680
rect 5128 38592 5136 38656
rect 5200 38592 5216 38656
rect 5280 38592 5296 38656
rect 5360 38592 5376 38656
rect 5440 38592 5448 38656
rect 5128 37568 5448 38592
rect 5128 37504 5136 37568
rect 5200 37504 5216 37568
rect 5280 37504 5296 37568
rect 5360 37504 5376 37568
rect 5440 37504 5448 37568
rect 5128 36480 5448 37504
rect 5128 36416 5136 36480
rect 5200 36416 5216 36480
rect 5280 36416 5296 36480
rect 5360 36416 5376 36480
rect 5440 36416 5448 36480
rect 5128 36260 5448 36416
rect 5128 36024 5170 36260
rect 5406 36024 5448 36260
rect 5128 35392 5448 36024
rect 5128 35328 5136 35392
rect 5200 35328 5216 35392
rect 5280 35328 5296 35392
rect 5360 35328 5376 35392
rect 5440 35328 5448 35392
rect 5128 34304 5448 35328
rect 5128 34240 5136 34304
rect 5200 34240 5216 34304
rect 5280 34240 5296 34304
rect 5360 34240 5376 34304
rect 5440 34240 5448 34304
rect 5128 33216 5448 34240
rect 5128 33152 5136 33216
rect 5200 33152 5216 33216
rect 5280 33152 5296 33216
rect 5360 33152 5376 33216
rect 5440 33152 5448 33216
rect 5128 32128 5448 33152
rect 5128 32064 5136 32128
rect 5200 32064 5216 32128
rect 5280 32064 5296 32128
rect 5360 32064 5376 32128
rect 5440 32064 5448 32128
rect 5128 31040 5448 32064
rect 5128 30976 5136 31040
rect 5200 30976 5216 31040
rect 5280 30976 5296 31040
rect 5360 30976 5376 31040
rect 5440 30976 5448 31040
rect 5128 29952 5448 30976
rect 5128 29888 5136 29952
rect 5200 29888 5216 29952
rect 5280 29888 5296 29952
rect 5360 29888 5376 29952
rect 5440 29888 5448 29952
rect 5128 28864 5448 29888
rect 5128 28800 5136 28864
rect 5200 28800 5216 28864
rect 5280 28800 5296 28864
rect 5360 28800 5376 28864
rect 5440 28800 5448 28864
rect 5128 27776 5448 28800
rect 5128 27712 5136 27776
rect 5200 27712 5216 27776
rect 5280 27712 5296 27776
rect 5360 27712 5376 27776
rect 5440 27712 5448 27776
rect 5128 26688 5448 27712
rect 5128 26624 5136 26688
rect 5200 26624 5216 26688
rect 5280 26624 5296 26688
rect 5360 26624 5376 26688
rect 5440 26624 5448 26688
rect 5128 25600 5448 26624
rect 5128 25536 5136 25600
rect 5200 25536 5216 25600
rect 5280 25536 5296 25600
rect 5360 25536 5376 25600
rect 5440 25536 5448 25600
rect 5128 24512 5448 25536
rect 5128 24448 5136 24512
rect 5200 24448 5216 24512
rect 5280 24448 5296 24512
rect 5360 24448 5376 24512
rect 5440 24448 5448 24512
rect 5128 23424 5448 24448
rect 5128 23360 5136 23424
rect 5200 23360 5216 23424
rect 5280 23360 5296 23424
rect 5360 23360 5376 23424
rect 5440 23360 5448 23424
rect 5128 22336 5448 23360
rect 5128 22272 5136 22336
rect 5200 22272 5216 22336
rect 5280 22272 5296 22336
rect 5360 22272 5376 22336
rect 5440 22272 5448 22336
rect 5128 21248 5448 22272
rect 5128 21184 5136 21248
rect 5200 21184 5216 21248
rect 5280 21184 5296 21248
rect 5360 21184 5376 21248
rect 5440 21184 5448 21248
rect 5128 20160 5448 21184
rect 5128 20096 5136 20160
rect 5200 20096 5216 20160
rect 5280 20096 5296 20160
rect 5360 20096 5376 20160
rect 5440 20096 5448 20160
rect 5128 19072 5448 20096
rect 5128 19008 5136 19072
rect 5200 19008 5216 19072
rect 5280 19008 5296 19072
rect 5360 19008 5376 19072
rect 5440 19008 5448 19072
rect 5128 17984 5448 19008
rect 5128 17920 5136 17984
rect 5200 17920 5216 17984
rect 5280 17920 5296 17984
rect 5360 17920 5376 17984
rect 5440 17920 5448 17984
rect 5128 16896 5448 17920
rect 5128 16832 5136 16896
rect 5200 16832 5216 16896
rect 5280 16832 5296 16896
rect 5360 16832 5376 16896
rect 5440 16832 5448 16896
rect 5128 15808 5448 16832
rect 5128 15744 5136 15808
rect 5200 15744 5216 15808
rect 5280 15744 5296 15808
rect 5360 15744 5376 15808
rect 5440 15744 5448 15808
rect 5128 14720 5448 15744
rect 5128 14656 5136 14720
rect 5200 14656 5216 14720
rect 5280 14656 5296 14720
rect 5360 14656 5376 14720
rect 5440 14656 5448 14720
rect 5128 13632 5448 14656
rect 5128 13568 5136 13632
rect 5200 13568 5216 13632
rect 5280 13568 5296 13632
rect 5360 13568 5376 13632
rect 5440 13568 5448 13632
rect 5128 12544 5448 13568
rect 5128 12480 5136 12544
rect 5200 12480 5216 12544
rect 5280 12480 5296 12544
rect 5360 12480 5376 12544
rect 5440 12480 5448 12544
rect 5128 11456 5448 12480
rect 5128 11392 5136 11456
rect 5200 11392 5216 11456
rect 5280 11392 5296 11456
rect 5360 11392 5376 11456
rect 5440 11392 5448 11456
rect 5128 10368 5448 11392
rect 5128 10304 5136 10368
rect 5200 10304 5216 10368
rect 5280 10304 5296 10368
rect 5360 10304 5376 10368
rect 5440 10304 5448 10368
rect 5128 9280 5448 10304
rect 5128 9216 5136 9280
rect 5200 9216 5216 9280
rect 5280 9216 5296 9280
rect 5360 9216 5376 9280
rect 5440 9216 5448 9280
rect 5128 8192 5448 9216
rect 5128 8128 5136 8192
rect 5200 8128 5216 8192
rect 5280 8128 5296 8192
rect 5360 8128 5376 8192
rect 5440 8128 5448 8192
rect 5128 7104 5448 8128
rect 5128 7040 5136 7104
rect 5200 7040 5216 7104
rect 5280 7040 5296 7104
rect 5360 7040 5376 7104
rect 5440 7040 5448 7104
rect 5128 6016 5448 7040
rect 5128 5952 5136 6016
rect 5200 5952 5216 6016
rect 5280 5952 5296 6016
rect 5360 5952 5376 6016
rect 5440 5952 5448 6016
rect 5128 5624 5448 5952
rect 5128 5388 5170 5624
rect 5406 5388 5448 5624
rect 5128 4928 5448 5388
rect 5128 4864 5136 4928
rect 5200 4864 5216 4928
rect 5280 4864 5296 4928
rect 5360 4864 5376 4928
rect 5440 4864 5448 4928
rect 5128 3840 5448 4864
rect 5128 3776 5136 3840
rect 5200 3776 5216 3840
rect 5280 3776 5296 3840
rect 5360 3776 5376 3840
rect 5440 3776 5448 3840
rect 5128 2752 5448 3776
rect 5128 2688 5136 2752
rect 5200 2688 5216 2752
rect 5280 2688 5296 2752
rect 5360 2688 5376 2752
rect 5440 2688 5448 2752
rect 5128 2128 5448 2688
rect 5788 77280 6108 77840
rect 5788 77216 5796 77280
rect 5860 77216 5876 77280
rect 5940 77216 5956 77280
rect 6020 77216 6036 77280
rect 6100 77216 6108 77280
rect 5788 76192 6108 77216
rect 5788 76128 5796 76192
rect 5860 76128 5876 76192
rect 5940 76128 5956 76192
rect 6020 76128 6036 76192
rect 6100 76128 6108 76192
rect 5788 75104 6108 76128
rect 5788 75040 5796 75104
rect 5860 75040 5876 75104
rect 5940 75040 5956 75104
rect 6020 75040 6036 75104
rect 6100 75040 6108 75104
rect 5788 74016 6108 75040
rect 5788 73952 5796 74016
rect 5860 73952 5876 74016
rect 5940 73952 5956 74016
rect 6020 73952 6036 74016
rect 6100 73952 6108 74016
rect 5788 72928 6108 73952
rect 5788 72864 5796 72928
rect 5860 72864 5876 72928
rect 5940 72864 5956 72928
rect 6020 72864 6036 72928
rect 6100 72864 6108 72928
rect 5788 71840 6108 72864
rect 5788 71776 5796 71840
rect 5860 71776 5876 71840
rect 5940 71776 5956 71840
rect 6020 71776 6036 71840
rect 6100 71776 6108 71840
rect 5788 70752 6108 71776
rect 5788 70688 5796 70752
rect 5860 70688 5876 70752
rect 5940 70688 5956 70752
rect 6020 70688 6036 70752
rect 6100 70688 6108 70752
rect 5788 69664 6108 70688
rect 5788 69600 5796 69664
rect 5860 69600 5876 69664
rect 5940 69600 5956 69664
rect 6020 69600 6036 69664
rect 6100 69600 6108 69664
rect 5788 68576 6108 69600
rect 5788 68512 5796 68576
rect 5860 68512 5876 68576
rect 5940 68512 5956 68576
rect 6020 68512 6036 68576
rect 6100 68512 6108 68576
rect 5788 67556 6108 68512
rect 5788 67488 5830 67556
rect 6066 67488 6108 67556
rect 5788 67424 5796 67488
rect 6100 67424 6108 67488
rect 5788 67320 5830 67424
rect 6066 67320 6108 67424
rect 5788 66400 6108 67320
rect 5788 66336 5796 66400
rect 5860 66336 5876 66400
rect 5940 66336 5956 66400
rect 6020 66336 6036 66400
rect 6100 66336 6108 66400
rect 5788 65312 6108 66336
rect 5788 65248 5796 65312
rect 5860 65248 5876 65312
rect 5940 65248 5956 65312
rect 6020 65248 6036 65312
rect 6100 65248 6108 65312
rect 5788 64224 6108 65248
rect 5788 64160 5796 64224
rect 5860 64160 5876 64224
rect 5940 64160 5956 64224
rect 6020 64160 6036 64224
rect 6100 64160 6108 64224
rect 5788 63136 6108 64160
rect 5788 63072 5796 63136
rect 5860 63072 5876 63136
rect 5940 63072 5956 63136
rect 6020 63072 6036 63136
rect 6100 63072 6108 63136
rect 5788 62048 6108 63072
rect 5788 61984 5796 62048
rect 5860 61984 5876 62048
rect 5940 61984 5956 62048
rect 6020 61984 6036 62048
rect 6100 61984 6108 62048
rect 5788 60960 6108 61984
rect 5788 60896 5796 60960
rect 5860 60896 5876 60960
rect 5940 60896 5956 60960
rect 6020 60896 6036 60960
rect 6100 60896 6108 60960
rect 5788 59872 6108 60896
rect 5788 59808 5796 59872
rect 5860 59808 5876 59872
rect 5940 59808 5956 59872
rect 6020 59808 6036 59872
rect 6100 59808 6108 59872
rect 5788 58784 6108 59808
rect 5788 58720 5796 58784
rect 5860 58720 5876 58784
rect 5940 58720 5956 58784
rect 6020 58720 6036 58784
rect 6100 58720 6108 58784
rect 5788 57696 6108 58720
rect 5788 57632 5796 57696
rect 5860 57632 5876 57696
rect 5940 57632 5956 57696
rect 6020 57632 6036 57696
rect 6100 57632 6108 57696
rect 5788 56608 6108 57632
rect 5788 56544 5796 56608
rect 5860 56544 5876 56608
rect 5940 56544 5956 56608
rect 6020 56544 6036 56608
rect 6100 56544 6108 56608
rect 5788 55520 6108 56544
rect 5788 55456 5796 55520
rect 5860 55456 5876 55520
rect 5940 55456 5956 55520
rect 6020 55456 6036 55520
rect 6100 55456 6108 55520
rect 5788 54432 6108 55456
rect 5788 54368 5796 54432
rect 5860 54368 5876 54432
rect 5940 54368 5956 54432
rect 6020 54368 6036 54432
rect 6100 54368 6108 54432
rect 5788 53344 6108 54368
rect 5788 53280 5796 53344
rect 5860 53280 5876 53344
rect 5940 53280 5956 53344
rect 6020 53280 6036 53344
rect 6100 53280 6108 53344
rect 5788 52256 6108 53280
rect 5788 52192 5796 52256
rect 5860 52192 5876 52256
rect 5940 52192 5956 52256
rect 6020 52192 6036 52256
rect 6100 52192 6108 52256
rect 5788 51168 6108 52192
rect 5788 51104 5796 51168
rect 5860 51104 5876 51168
rect 5940 51104 5956 51168
rect 6020 51104 6036 51168
rect 6100 51104 6108 51168
rect 5788 50080 6108 51104
rect 5788 50016 5796 50080
rect 5860 50016 5876 50080
rect 5940 50016 5956 50080
rect 6020 50016 6036 50080
rect 6100 50016 6108 50080
rect 5788 48992 6108 50016
rect 5788 48928 5796 48992
rect 5860 48928 5876 48992
rect 5940 48928 5956 48992
rect 6020 48928 6036 48992
rect 6100 48928 6108 48992
rect 5788 47904 6108 48928
rect 5788 47840 5796 47904
rect 5860 47840 5876 47904
rect 5940 47840 5956 47904
rect 6020 47840 6036 47904
rect 6100 47840 6108 47904
rect 5788 46816 6108 47840
rect 5788 46752 5796 46816
rect 5860 46752 5876 46816
rect 5940 46752 5956 46816
rect 6020 46752 6036 46816
rect 6100 46752 6108 46816
rect 5788 45728 6108 46752
rect 5788 45664 5796 45728
rect 5860 45664 5876 45728
rect 5940 45664 5956 45728
rect 6020 45664 6036 45728
rect 6100 45664 6108 45728
rect 5788 44640 6108 45664
rect 5788 44576 5796 44640
rect 5860 44576 5876 44640
rect 5940 44576 5956 44640
rect 6020 44576 6036 44640
rect 6100 44576 6108 44640
rect 5788 43552 6108 44576
rect 5788 43488 5796 43552
rect 5860 43488 5876 43552
rect 5940 43488 5956 43552
rect 6020 43488 6036 43552
rect 6100 43488 6108 43552
rect 5788 42464 6108 43488
rect 5788 42400 5796 42464
rect 5860 42400 5876 42464
rect 5940 42400 5956 42464
rect 6020 42400 6036 42464
rect 6100 42400 6108 42464
rect 5788 41376 6108 42400
rect 5788 41312 5796 41376
rect 5860 41312 5876 41376
rect 5940 41312 5956 41376
rect 6020 41312 6036 41376
rect 6100 41312 6108 41376
rect 5788 40288 6108 41312
rect 5788 40224 5796 40288
rect 5860 40224 5876 40288
rect 5940 40224 5956 40288
rect 6020 40224 6036 40288
rect 6100 40224 6108 40288
rect 5788 39200 6108 40224
rect 5788 39136 5796 39200
rect 5860 39136 5876 39200
rect 5940 39136 5956 39200
rect 6020 39136 6036 39200
rect 6100 39136 6108 39200
rect 5788 38112 6108 39136
rect 5788 38048 5796 38112
rect 5860 38048 5876 38112
rect 5940 38048 5956 38112
rect 6020 38048 6036 38112
rect 6100 38048 6108 38112
rect 5788 37024 6108 38048
rect 5788 36960 5796 37024
rect 5860 36960 5876 37024
rect 5940 36960 5956 37024
rect 6020 36960 6036 37024
rect 6100 36960 6108 37024
rect 5788 36920 6108 36960
rect 5788 36684 5830 36920
rect 6066 36684 6108 36920
rect 5788 35936 6108 36684
rect 5788 35872 5796 35936
rect 5860 35872 5876 35936
rect 5940 35872 5956 35936
rect 6020 35872 6036 35936
rect 6100 35872 6108 35936
rect 5788 34848 6108 35872
rect 5788 34784 5796 34848
rect 5860 34784 5876 34848
rect 5940 34784 5956 34848
rect 6020 34784 6036 34848
rect 6100 34784 6108 34848
rect 5788 33760 6108 34784
rect 5788 33696 5796 33760
rect 5860 33696 5876 33760
rect 5940 33696 5956 33760
rect 6020 33696 6036 33760
rect 6100 33696 6108 33760
rect 5788 32672 6108 33696
rect 5788 32608 5796 32672
rect 5860 32608 5876 32672
rect 5940 32608 5956 32672
rect 6020 32608 6036 32672
rect 6100 32608 6108 32672
rect 5788 31584 6108 32608
rect 5788 31520 5796 31584
rect 5860 31520 5876 31584
rect 5940 31520 5956 31584
rect 6020 31520 6036 31584
rect 6100 31520 6108 31584
rect 5788 30496 6108 31520
rect 5788 30432 5796 30496
rect 5860 30432 5876 30496
rect 5940 30432 5956 30496
rect 6020 30432 6036 30496
rect 6100 30432 6108 30496
rect 5788 29408 6108 30432
rect 5788 29344 5796 29408
rect 5860 29344 5876 29408
rect 5940 29344 5956 29408
rect 6020 29344 6036 29408
rect 6100 29344 6108 29408
rect 5788 28320 6108 29344
rect 5788 28256 5796 28320
rect 5860 28256 5876 28320
rect 5940 28256 5956 28320
rect 6020 28256 6036 28320
rect 6100 28256 6108 28320
rect 5788 27232 6108 28256
rect 5788 27168 5796 27232
rect 5860 27168 5876 27232
rect 5940 27168 5956 27232
rect 6020 27168 6036 27232
rect 6100 27168 6108 27232
rect 5788 26144 6108 27168
rect 5788 26080 5796 26144
rect 5860 26080 5876 26144
rect 5940 26080 5956 26144
rect 6020 26080 6036 26144
rect 6100 26080 6108 26144
rect 5788 25056 6108 26080
rect 5788 24992 5796 25056
rect 5860 24992 5876 25056
rect 5940 24992 5956 25056
rect 6020 24992 6036 25056
rect 6100 24992 6108 25056
rect 5788 23968 6108 24992
rect 5788 23904 5796 23968
rect 5860 23904 5876 23968
rect 5940 23904 5956 23968
rect 6020 23904 6036 23968
rect 6100 23904 6108 23968
rect 5788 22880 6108 23904
rect 5788 22816 5796 22880
rect 5860 22816 5876 22880
rect 5940 22816 5956 22880
rect 6020 22816 6036 22880
rect 6100 22816 6108 22880
rect 5788 21792 6108 22816
rect 5788 21728 5796 21792
rect 5860 21728 5876 21792
rect 5940 21728 5956 21792
rect 6020 21728 6036 21792
rect 6100 21728 6108 21792
rect 5788 20704 6108 21728
rect 5788 20640 5796 20704
rect 5860 20640 5876 20704
rect 5940 20640 5956 20704
rect 6020 20640 6036 20704
rect 6100 20640 6108 20704
rect 5788 19616 6108 20640
rect 5788 19552 5796 19616
rect 5860 19552 5876 19616
rect 5940 19552 5956 19616
rect 6020 19552 6036 19616
rect 6100 19552 6108 19616
rect 5788 18528 6108 19552
rect 5788 18464 5796 18528
rect 5860 18464 5876 18528
rect 5940 18464 5956 18528
rect 6020 18464 6036 18528
rect 6100 18464 6108 18528
rect 5788 17440 6108 18464
rect 5788 17376 5796 17440
rect 5860 17376 5876 17440
rect 5940 17376 5956 17440
rect 6020 17376 6036 17440
rect 6100 17376 6108 17440
rect 5788 16352 6108 17376
rect 5788 16288 5796 16352
rect 5860 16288 5876 16352
rect 5940 16288 5956 16352
rect 6020 16288 6036 16352
rect 6100 16288 6108 16352
rect 5788 15264 6108 16288
rect 5788 15200 5796 15264
rect 5860 15200 5876 15264
rect 5940 15200 5956 15264
rect 6020 15200 6036 15264
rect 6100 15200 6108 15264
rect 5788 14176 6108 15200
rect 5788 14112 5796 14176
rect 5860 14112 5876 14176
rect 5940 14112 5956 14176
rect 6020 14112 6036 14176
rect 6100 14112 6108 14176
rect 5788 13088 6108 14112
rect 5788 13024 5796 13088
rect 5860 13024 5876 13088
rect 5940 13024 5956 13088
rect 6020 13024 6036 13088
rect 6100 13024 6108 13088
rect 5788 12000 6108 13024
rect 5788 11936 5796 12000
rect 5860 11936 5876 12000
rect 5940 11936 5956 12000
rect 6020 11936 6036 12000
rect 6100 11936 6108 12000
rect 5788 10912 6108 11936
rect 5788 10848 5796 10912
rect 5860 10848 5876 10912
rect 5940 10848 5956 10912
rect 6020 10848 6036 10912
rect 6100 10848 6108 10912
rect 5788 9824 6108 10848
rect 5788 9760 5796 9824
rect 5860 9760 5876 9824
rect 5940 9760 5956 9824
rect 6020 9760 6036 9824
rect 6100 9760 6108 9824
rect 5788 8736 6108 9760
rect 5788 8672 5796 8736
rect 5860 8672 5876 8736
rect 5940 8672 5956 8736
rect 6020 8672 6036 8736
rect 6100 8672 6108 8736
rect 5788 7648 6108 8672
rect 5788 7584 5796 7648
rect 5860 7584 5876 7648
rect 5940 7584 5956 7648
rect 6020 7584 6036 7648
rect 6100 7584 6108 7648
rect 5788 6560 6108 7584
rect 5788 6496 5796 6560
rect 5860 6496 5876 6560
rect 5940 6496 5956 6560
rect 6020 6496 6036 6560
rect 6100 6496 6108 6560
rect 5788 6284 6108 6496
rect 5788 6048 5830 6284
rect 6066 6048 6108 6284
rect 5788 5472 6108 6048
rect 5788 5408 5796 5472
rect 5860 5408 5876 5472
rect 5940 5408 5956 5472
rect 6020 5408 6036 5472
rect 6100 5408 6108 5472
rect 5788 4384 6108 5408
rect 5788 4320 5796 4384
rect 5860 4320 5876 4384
rect 5940 4320 5956 4384
rect 6020 4320 6036 4384
rect 6100 4320 6108 4384
rect 5788 3296 6108 4320
rect 5788 3232 5796 3296
rect 5860 3232 5876 3296
rect 5940 3232 5956 3296
rect 6020 3232 6036 3296
rect 6100 3232 6108 3296
rect 5788 2208 6108 3232
rect 5788 2144 5796 2208
rect 5860 2144 5876 2208
rect 5940 2144 5956 2208
rect 6020 2144 6036 2208
rect 6100 2144 6108 2208
rect 5788 2128 6108 2144
rect 35848 77824 36168 77840
rect 35848 77760 35856 77824
rect 35920 77760 35936 77824
rect 36000 77760 36016 77824
rect 36080 77760 36096 77824
rect 36160 77760 36168 77824
rect 35848 76736 36168 77760
rect 35848 76672 35856 76736
rect 35920 76672 35936 76736
rect 36000 76672 36016 76736
rect 36080 76672 36096 76736
rect 36160 76672 36168 76736
rect 35848 75648 36168 76672
rect 35848 75584 35856 75648
rect 35920 75584 35936 75648
rect 36000 75584 36016 75648
rect 36080 75584 36096 75648
rect 36160 75584 36168 75648
rect 35848 74560 36168 75584
rect 35848 74496 35856 74560
rect 35920 74496 35936 74560
rect 36000 74496 36016 74560
rect 36080 74496 36096 74560
rect 36160 74496 36168 74560
rect 35848 73472 36168 74496
rect 35848 73408 35856 73472
rect 35920 73408 35936 73472
rect 36000 73408 36016 73472
rect 36080 73408 36096 73472
rect 36160 73408 36168 73472
rect 35848 72384 36168 73408
rect 35848 72320 35856 72384
rect 35920 72320 35936 72384
rect 36000 72320 36016 72384
rect 36080 72320 36096 72384
rect 36160 72320 36168 72384
rect 35848 71296 36168 72320
rect 35848 71232 35856 71296
rect 35920 71232 35936 71296
rect 36000 71232 36016 71296
rect 36080 71232 36096 71296
rect 36160 71232 36168 71296
rect 35848 70208 36168 71232
rect 35848 70144 35856 70208
rect 35920 70144 35936 70208
rect 36000 70144 36016 70208
rect 36080 70144 36096 70208
rect 36160 70144 36168 70208
rect 35848 69120 36168 70144
rect 35848 69056 35856 69120
rect 35920 69056 35936 69120
rect 36000 69056 36016 69120
rect 36080 69056 36096 69120
rect 36160 69056 36168 69120
rect 35848 68032 36168 69056
rect 35848 67968 35856 68032
rect 35920 67968 35936 68032
rect 36000 67968 36016 68032
rect 36080 67968 36096 68032
rect 36160 67968 36168 68032
rect 35848 66944 36168 67968
rect 35848 66880 35856 66944
rect 35920 66896 35936 66944
rect 36000 66896 36016 66944
rect 36080 66896 36096 66944
rect 36160 66880 36168 66944
rect 35848 66660 35890 66880
rect 36126 66660 36168 66880
rect 35848 65856 36168 66660
rect 35848 65792 35856 65856
rect 35920 65792 35936 65856
rect 36000 65792 36016 65856
rect 36080 65792 36096 65856
rect 36160 65792 36168 65856
rect 35848 64768 36168 65792
rect 35848 64704 35856 64768
rect 35920 64704 35936 64768
rect 36000 64704 36016 64768
rect 36080 64704 36096 64768
rect 36160 64704 36168 64768
rect 35848 63680 36168 64704
rect 35848 63616 35856 63680
rect 35920 63616 35936 63680
rect 36000 63616 36016 63680
rect 36080 63616 36096 63680
rect 36160 63616 36168 63680
rect 35848 62592 36168 63616
rect 35848 62528 35856 62592
rect 35920 62528 35936 62592
rect 36000 62528 36016 62592
rect 36080 62528 36096 62592
rect 36160 62528 36168 62592
rect 35848 61504 36168 62528
rect 35848 61440 35856 61504
rect 35920 61440 35936 61504
rect 36000 61440 36016 61504
rect 36080 61440 36096 61504
rect 36160 61440 36168 61504
rect 35848 60416 36168 61440
rect 35848 60352 35856 60416
rect 35920 60352 35936 60416
rect 36000 60352 36016 60416
rect 36080 60352 36096 60416
rect 36160 60352 36168 60416
rect 35848 59328 36168 60352
rect 35848 59264 35856 59328
rect 35920 59264 35936 59328
rect 36000 59264 36016 59328
rect 36080 59264 36096 59328
rect 36160 59264 36168 59328
rect 35848 58240 36168 59264
rect 35848 58176 35856 58240
rect 35920 58176 35936 58240
rect 36000 58176 36016 58240
rect 36080 58176 36096 58240
rect 36160 58176 36168 58240
rect 35848 57152 36168 58176
rect 35848 57088 35856 57152
rect 35920 57088 35936 57152
rect 36000 57088 36016 57152
rect 36080 57088 36096 57152
rect 36160 57088 36168 57152
rect 35848 56064 36168 57088
rect 35848 56000 35856 56064
rect 35920 56000 35936 56064
rect 36000 56000 36016 56064
rect 36080 56000 36096 56064
rect 36160 56000 36168 56064
rect 35848 54976 36168 56000
rect 35848 54912 35856 54976
rect 35920 54912 35936 54976
rect 36000 54912 36016 54976
rect 36080 54912 36096 54976
rect 36160 54912 36168 54976
rect 35848 53888 36168 54912
rect 35848 53824 35856 53888
rect 35920 53824 35936 53888
rect 36000 53824 36016 53888
rect 36080 53824 36096 53888
rect 36160 53824 36168 53888
rect 35848 52800 36168 53824
rect 35848 52736 35856 52800
rect 35920 52736 35936 52800
rect 36000 52736 36016 52800
rect 36080 52736 36096 52800
rect 36160 52736 36168 52800
rect 35848 51712 36168 52736
rect 35848 51648 35856 51712
rect 35920 51648 35936 51712
rect 36000 51648 36016 51712
rect 36080 51648 36096 51712
rect 36160 51648 36168 51712
rect 35848 50624 36168 51648
rect 35848 50560 35856 50624
rect 35920 50560 35936 50624
rect 36000 50560 36016 50624
rect 36080 50560 36096 50624
rect 36160 50560 36168 50624
rect 35848 49536 36168 50560
rect 35848 49472 35856 49536
rect 35920 49472 35936 49536
rect 36000 49472 36016 49536
rect 36080 49472 36096 49536
rect 36160 49472 36168 49536
rect 35848 48448 36168 49472
rect 35848 48384 35856 48448
rect 35920 48384 35936 48448
rect 36000 48384 36016 48448
rect 36080 48384 36096 48448
rect 36160 48384 36168 48448
rect 35848 47360 36168 48384
rect 35848 47296 35856 47360
rect 35920 47296 35936 47360
rect 36000 47296 36016 47360
rect 36080 47296 36096 47360
rect 36160 47296 36168 47360
rect 35848 46272 36168 47296
rect 35848 46208 35856 46272
rect 35920 46208 35936 46272
rect 36000 46208 36016 46272
rect 36080 46208 36096 46272
rect 36160 46208 36168 46272
rect 35848 45184 36168 46208
rect 35848 45120 35856 45184
rect 35920 45120 35936 45184
rect 36000 45120 36016 45184
rect 36080 45120 36096 45184
rect 36160 45120 36168 45184
rect 35848 44096 36168 45120
rect 35848 44032 35856 44096
rect 35920 44032 35936 44096
rect 36000 44032 36016 44096
rect 36080 44032 36096 44096
rect 36160 44032 36168 44096
rect 35848 43008 36168 44032
rect 35848 42944 35856 43008
rect 35920 42944 35936 43008
rect 36000 42944 36016 43008
rect 36080 42944 36096 43008
rect 36160 42944 36168 43008
rect 35848 41920 36168 42944
rect 35848 41856 35856 41920
rect 35920 41856 35936 41920
rect 36000 41856 36016 41920
rect 36080 41856 36096 41920
rect 36160 41856 36168 41920
rect 35848 40832 36168 41856
rect 35848 40768 35856 40832
rect 35920 40768 35936 40832
rect 36000 40768 36016 40832
rect 36080 40768 36096 40832
rect 36160 40768 36168 40832
rect 35848 39744 36168 40768
rect 35848 39680 35856 39744
rect 35920 39680 35936 39744
rect 36000 39680 36016 39744
rect 36080 39680 36096 39744
rect 36160 39680 36168 39744
rect 35848 38656 36168 39680
rect 35848 38592 35856 38656
rect 35920 38592 35936 38656
rect 36000 38592 36016 38656
rect 36080 38592 36096 38656
rect 36160 38592 36168 38656
rect 35848 37568 36168 38592
rect 35848 37504 35856 37568
rect 35920 37504 35936 37568
rect 36000 37504 36016 37568
rect 36080 37504 36096 37568
rect 36160 37504 36168 37568
rect 35848 36480 36168 37504
rect 35848 36416 35856 36480
rect 35920 36416 35936 36480
rect 36000 36416 36016 36480
rect 36080 36416 36096 36480
rect 36160 36416 36168 36480
rect 35848 36260 36168 36416
rect 35848 36024 35890 36260
rect 36126 36024 36168 36260
rect 35848 35392 36168 36024
rect 35848 35328 35856 35392
rect 35920 35328 35936 35392
rect 36000 35328 36016 35392
rect 36080 35328 36096 35392
rect 36160 35328 36168 35392
rect 35848 34304 36168 35328
rect 35848 34240 35856 34304
rect 35920 34240 35936 34304
rect 36000 34240 36016 34304
rect 36080 34240 36096 34304
rect 36160 34240 36168 34304
rect 35848 33216 36168 34240
rect 35848 33152 35856 33216
rect 35920 33152 35936 33216
rect 36000 33152 36016 33216
rect 36080 33152 36096 33216
rect 36160 33152 36168 33216
rect 35848 32128 36168 33152
rect 35848 32064 35856 32128
rect 35920 32064 35936 32128
rect 36000 32064 36016 32128
rect 36080 32064 36096 32128
rect 36160 32064 36168 32128
rect 35848 31040 36168 32064
rect 35848 30976 35856 31040
rect 35920 30976 35936 31040
rect 36000 30976 36016 31040
rect 36080 30976 36096 31040
rect 36160 30976 36168 31040
rect 35848 29952 36168 30976
rect 35848 29888 35856 29952
rect 35920 29888 35936 29952
rect 36000 29888 36016 29952
rect 36080 29888 36096 29952
rect 36160 29888 36168 29952
rect 35848 28864 36168 29888
rect 35848 28800 35856 28864
rect 35920 28800 35936 28864
rect 36000 28800 36016 28864
rect 36080 28800 36096 28864
rect 36160 28800 36168 28864
rect 35848 27776 36168 28800
rect 35848 27712 35856 27776
rect 35920 27712 35936 27776
rect 36000 27712 36016 27776
rect 36080 27712 36096 27776
rect 36160 27712 36168 27776
rect 35848 26688 36168 27712
rect 35848 26624 35856 26688
rect 35920 26624 35936 26688
rect 36000 26624 36016 26688
rect 36080 26624 36096 26688
rect 36160 26624 36168 26688
rect 35848 25600 36168 26624
rect 35848 25536 35856 25600
rect 35920 25536 35936 25600
rect 36000 25536 36016 25600
rect 36080 25536 36096 25600
rect 36160 25536 36168 25600
rect 35848 24512 36168 25536
rect 35848 24448 35856 24512
rect 35920 24448 35936 24512
rect 36000 24448 36016 24512
rect 36080 24448 36096 24512
rect 36160 24448 36168 24512
rect 35848 23424 36168 24448
rect 35848 23360 35856 23424
rect 35920 23360 35936 23424
rect 36000 23360 36016 23424
rect 36080 23360 36096 23424
rect 36160 23360 36168 23424
rect 35848 22336 36168 23360
rect 35848 22272 35856 22336
rect 35920 22272 35936 22336
rect 36000 22272 36016 22336
rect 36080 22272 36096 22336
rect 36160 22272 36168 22336
rect 35848 21248 36168 22272
rect 35848 21184 35856 21248
rect 35920 21184 35936 21248
rect 36000 21184 36016 21248
rect 36080 21184 36096 21248
rect 36160 21184 36168 21248
rect 35848 20160 36168 21184
rect 35848 20096 35856 20160
rect 35920 20096 35936 20160
rect 36000 20096 36016 20160
rect 36080 20096 36096 20160
rect 36160 20096 36168 20160
rect 35848 19072 36168 20096
rect 35848 19008 35856 19072
rect 35920 19008 35936 19072
rect 36000 19008 36016 19072
rect 36080 19008 36096 19072
rect 36160 19008 36168 19072
rect 35848 17984 36168 19008
rect 35848 17920 35856 17984
rect 35920 17920 35936 17984
rect 36000 17920 36016 17984
rect 36080 17920 36096 17984
rect 36160 17920 36168 17984
rect 35848 16896 36168 17920
rect 35848 16832 35856 16896
rect 35920 16832 35936 16896
rect 36000 16832 36016 16896
rect 36080 16832 36096 16896
rect 36160 16832 36168 16896
rect 35848 15808 36168 16832
rect 35848 15744 35856 15808
rect 35920 15744 35936 15808
rect 36000 15744 36016 15808
rect 36080 15744 36096 15808
rect 36160 15744 36168 15808
rect 35848 14720 36168 15744
rect 35848 14656 35856 14720
rect 35920 14656 35936 14720
rect 36000 14656 36016 14720
rect 36080 14656 36096 14720
rect 36160 14656 36168 14720
rect 35848 13632 36168 14656
rect 35848 13568 35856 13632
rect 35920 13568 35936 13632
rect 36000 13568 36016 13632
rect 36080 13568 36096 13632
rect 36160 13568 36168 13632
rect 35848 12544 36168 13568
rect 35848 12480 35856 12544
rect 35920 12480 35936 12544
rect 36000 12480 36016 12544
rect 36080 12480 36096 12544
rect 36160 12480 36168 12544
rect 35848 11456 36168 12480
rect 35848 11392 35856 11456
rect 35920 11392 35936 11456
rect 36000 11392 36016 11456
rect 36080 11392 36096 11456
rect 36160 11392 36168 11456
rect 35848 10368 36168 11392
rect 35848 10304 35856 10368
rect 35920 10304 35936 10368
rect 36000 10304 36016 10368
rect 36080 10304 36096 10368
rect 36160 10304 36168 10368
rect 35848 9280 36168 10304
rect 35848 9216 35856 9280
rect 35920 9216 35936 9280
rect 36000 9216 36016 9280
rect 36080 9216 36096 9280
rect 36160 9216 36168 9280
rect 35848 8192 36168 9216
rect 35848 8128 35856 8192
rect 35920 8128 35936 8192
rect 36000 8128 36016 8192
rect 36080 8128 36096 8192
rect 36160 8128 36168 8192
rect 35848 7104 36168 8128
rect 35848 7040 35856 7104
rect 35920 7040 35936 7104
rect 36000 7040 36016 7104
rect 36080 7040 36096 7104
rect 36160 7040 36168 7104
rect 35848 6016 36168 7040
rect 35848 5952 35856 6016
rect 35920 5952 35936 6016
rect 36000 5952 36016 6016
rect 36080 5952 36096 6016
rect 36160 5952 36168 6016
rect 35848 5624 36168 5952
rect 35848 5388 35890 5624
rect 36126 5388 36168 5624
rect 35848 4928 36168 5388
rect 35848 4864 35856 4928
rect 35920 4864 35936 4928
rect 36000 4864 36016 4928
rect 36080 4864 36096 4928
rect 36160 4864 36168 4928
rect 35848 3840 36168 4864
rect 35848 3776 35856 3840
rect 35920 3776 35936 3840
rect 36000 3776 36016 3840
rect 36080 3776 36096 3840
rect 36160 3776 36168 3840
rect 35848 2752 36168 3776
rect 35848 2688 35856 2752
rect 35920 2688 35936 2752
rect 36000 2688 36016 2752
rect 36080 2688 36096 2752
rect 36160 2688 36168 2752
rect 35848 2128 36168 2688
rect 36508 77280 36828 77840
rect 36508 77216 36516 77280
rect 36580 77216 36596 77280
rect 36660 77216 36676 77280
rect 36740 77216 36756 77280
rect 36820 77216 36828 77280
rect 36508 76192 36828 77216
rect 36508 76128 36516 76192
rect 36580 76128 36596 76192
rect 36660 76128 36676 76192
rect 36740 76128 36756 76192
rect 36820 76128 36828 76192
rect 36508 75104 36828 76128
rect 36508 75040 36516 75104
rect 36580 75040 36596 75104
rect 36660 75040 36676 75104
rect 36740 75040 36756 75104
rect 36820 75040 36828 75104
rect 36508 74016 36828 75040
rect 36508 73952 36516 74016
rect 36580 73952 36596 74016
rect 36660 73952 36676 74016
rect 36740 73952 36756 74016
rect 36820 73952 36828 74016
rect 36508 72928 36828 73952
rect 36508 72864 36516 72928
rect 36580 72864 36596 72928
rect 36660 72864 36676 72928
rect 36740 72864 36756 72928
rect 36820 72864 36828 72928
rect 36508 71840 36828 72864
rect 36508 71776 36516 71840
rect 36580 71776 36596 71840
rect 36660 71776 36676 71840
rect 36740 71776 36756 71840
rect 36820 71776 36828 71840
rect 36508 70752 36828 71776
rect 36508 70688 36516 70752
rect 36580 70688 36596 70752
rect 36660 70688 36676 70752
rect 36740 70688 36756 70752
rect 36820 70688 36828 70752
rect 36508 69664 36828 70688
rect 36508 69600 36516 69664
rect 36580 69600 36596 69664
rect 36660 69600 36676 69664
rect 36740 69600 36756 69664
rect 36820 69600 36828 69664
rect 36508 68576 36828 69600
rect 36508 68512 36516 68576
rect 36580 68512 36596 68576
rect 36660 68512 36676 68576
rect 36740 68512 36756 68576
rect 36820 68512 36828 68576
rect 36508 67556 36828 68512
rect 36508 67488 36550 67556
rect 36786 67488 36828 67556
rect 36508 67424 36516 67488
rect 36820 67424 36828 67488
rect 36508 67320 36550 67424
rect 36786 67320 36828 67424
rect 36508 66400 36828 67320
rect 36508 66336 36516 66400
rect 36580 66336 36596 66400
rect 36660 66336 36676 66400
rect 36740 66336 36756 66400
rect 36820 66336 36828 66400
rect 36508 65312 36828 66336
rect 36508 65248 36516 65312
rect 36580 65248 36596 65312
rect 36660 65248 36676 65312
rect 36740 65248 36756 65312
rect 36820 65248 36828 65312
rect 36508 64224 36828 65248
rect 36508 64160 36516 64224
rect 36580 64160 36596 64224
rect 36660 64160 36676 64224
rect 36740 64160 36756 64224
rect 36820 64160 36828 64224
rect 36508 63136 36828 64160
rect 36508 63072 36516 63136
rect 36580 63072 36596 63136
rect 36660 63072 36676 63136
rect 36740 63072 36756 63136
rect 36820 63072 36828 63136
rect 36508 62048 36828 63072
rect 36508 61984 36516 62048
rect 36580 61984 36596 62048
rect 36660 61984 36676 62048
rect 36740 61984 36756 62048
rect 36820 61984 36828 62048
rect 36508 60960 36828 61984
rect 36508 60896 36516 60960
rect 36580 60896 36596 60960
rect 36660 60896 36676 60960
rect 36740 60896 36756 60960
rect 36820 60896 36828 60960
rect 36508 59872 36828 60896
rect 36508 59808 36516 59872
rect 36580 59808 36596 59872
rect 36660 59808 36676 59872
rect 36740 59808 36756 59872
rect 36820 59808 36828 59872
rect 36508 58784 36828 59808
rect 36508 58720 36516 58784
rect 36580 58720 36596 58784
rect 36660 58720 36676 58784
rect 36740 58720 36756 58784
rect 36820 58720 36828 58784
rect 36508 57696 36828 58720
rect 36508 57632 36516 57696
rect 36580 57632 36596 57696
rect 36660 57632 36676 57696
rect 36740 57632 36756 57696
rect 36820 57632 36828 57696
rect 36508 56608 36828 57632
rect 36508 56544 36516 56608
rect 36580 56544 36596 56608
rect 36660 56544 36676 56608
rect 36740 56544 36756 56608
rect 36820 56544 36828 56608
rect 36508 55520 36828 56544
rect 36508 55456 36516 55520
rect 36580 55456 36596 55520
rect 36660 55456 36676 55520
rect 36740 55456 36756 55520
rect 36820 55456 36828 55520
rect 36508 54432 36828 55456
rect 36508 54368 36516 54432
rect 36580 54368 36596 54432
rect 36660 54368 36676 54432
rect 36740 54368 36756 54432
rect 36820 54368 36828 54432
rect 36508 53344 36828 54368
rect 36508 53280 36516 53344
rect 36580 53280 36596 53344
rect 36660 53280 36676 53344
rect 36740 53280 36756 53344
rect 36820 53280 36828 53344
rect 36508 52256 36828 53280
rect 36508 52192 36516 52256
rect 36580 52192 36596 52256
rect 36660 52192 36676 52256
rect 36740 52192 36756 52256
rect 36820 52192 36828 52256
rect 36508 51168 36828 52192
rect 36508 51104 36516 51168
rect 36580 51104 36596 51168
rect 36660 51104 36676 51168
rect 36740 51104 36756 51168
rect 36820 51104 36828 51168
rect 36508 50080 36828 51104
rect 36508 50016 36516 50080
rect 36580 50016 36596 50080
rect 36660 50016 36676 50080
rect 36740 50016 36756 50080
rect 36820 50016 36828 50080
rect 36508 48992 36828 50016
rect 36508 48928 36516 48992
rect 36580 48928 36596 48992
rect 36660 48928 36676 48992
rect 36740 48928 36756 48992
rect 36820 48928 36828 48992
rect 36508 47904 36828 48928
rect 36508 47840 36516 47904
rect 36580 47840 36596 47904
rect 36660 47840 36676 47904
rect 36740 47840 36756 47904
rect 36820 47840 36828 47904
rect 36508 46816 36828 47840
rect 36508 46752 36516 46816
rect 36580 46752 36596 46816
rect 36660 46752 36676 46816
rect 36740 46752 36756 46816
rect 36820 46752 36828 46816
rect 36508 45728 36828 46752
rect 36508 45664 36516 45728
rect 36580 45664 36596 45728
rect 36660 45664 36676 45728
rect 36740 45664 36756 45728
rect 36820 45664 36828 45728
rect 36508 44640 36828 45664
rect 36508 44576 36516 44640
rect 36580 44576 36596 44640
rect 36660 44576 36676 44640
rect 36740 44576 36756 44640
rect 36820 44576 36828 44640
rect 36508 43552 36828 44576
rect 36508 43488 36516 43552
rect 36580 43488 36596 43552
rect 36660 43488 36676 43552
rect 36740 43488 36756 43552
rect 36820 43488 36828 43552
rect 36508 42464 36828 43488
rect 36508 42400 36516 42464
rect 36580 42400 36596 42464
rect 36660 42400 36676 42464
rect 36740 42400 36756 42464
rect 36820 42400 36828 42464
rect 36508 41376 36828 42400
rect 36508 41312 36516 41376
rect 36580 41312 36596 41376
rect 36660 41312 36676 41376
rect 36740 41312 36756 41376
rect 36820 41312 36828 41376
rect 36508 40288 36828 41312
rect 36508 40224 36516 40288
rect 36580 40224 36596 40288
rect 36660 40224 36676 40288
rect 36740 40224 36756 40288
rect 36820 40224 36828 40288
rect 36508 39200 36828 40224
rect 36508 39136 36516 39200
rect 36580 39136 36596 39200
rect 36660 39136 36676 39200
rect 36740 39136 36756 39200
rect 36820 39136 36828 39200
rect 36508 38112 36828 39136
rect 36508 38048 36516 38112
rect 36580 38048 36596 38112
rect 36660 38048 36676 38112
rect 36740 38048 36756 38112
rect 36820 38048 36828 38112
rect 36508 37024 36828 38048
rect 36508 36960 36516 37024
rect 36580 36960 36596 37024
rect 36660 36960 36676 37024
rect 36740 36960 36756 37024
rect 36820 36960 36828 37024
rect 36508 36920 36828 36960
rect 36508 36684 36550 36920
rect 36786 36684 36828 36920
rect 36508 35936 36828 36684
rect 36508 35872 36516 35936
rect 36580 35872 36596 35936
rect 36660 35872 36676 35936
rect 36740 35872 36756 35936
rect 36820 35872 36828 35936
rect 36508 34848 36828 35872
rect 36508 34784 36516 34848
rect 36580 34784 36596 34848
rect 36660 34784 36676 34848
rect 36740 34784 36756 34848
rect 36820 34784 36828 34848
rect 36508 33760 36828 34784
rect 36508 33696 36516 33760
rect 36580 33696 36596 33760
rect 36660 33696 36676 33760
rect 36740 33696 36756 33760
rect 36820 33696 36828 33760
rect 36508 32672 36828 33696
rect 36508 32608 36516 32672
rect 36580 32608 36596 32672
rect 36660 32608 36676 32672
rect 36740 32608 36756 32672
rect 36820 32608 36828 32672
rect 36508 31584 36828 32608
rect 36508 31520 36516 31584
rect 36580 31520 36596 31584
rect 36660 31520 36676 31584
rect 36740 31520 36756 31584
rect 36820 31520 36828 31584
rect 36508 30496 36828 31520
rect 36508 30432 36516 30496
rect 36580 30432 36596 30496
rect 36660 30432 36676 30496
rect 36740 30432 36756 30496
rect 36820 30432 36828 30496
rect 36508 29408 36828 30432
rect 36508 29344 36516 29408
rect 36580 29344 36596 29408
rect 36660 29344 36676 29408
rect 36740 29344 36756 29408
rect 36820 29344 36828 29408
rect 36508 28320 36828 29344
rect 36508 28256 36516 28320
rect 36580 28256 36596 28320
rect 36660 28256 36676 28320
rect 36740 28256 36756 28320
rect 36820 28256 36828 28320
rect 36508 27232 36828 28256
rect 36508 27168 36516 27232
rect 36580 27168 36596 27232
rect 36660 27168 36676 27232
rect 36740 27168 36756 27232
rect 36820 27168 36828 27232
rect 36508 26144 36828 27168
rect 36508 26080 36516 26144
rect 36580 26080 36596 26144
rect 36660 26080 36676 26144
rect 36740 26080 36756 26144
rect 36820 26080 36828 26144
rect 36508 25056 36828 26080
rect 36508 24992 36516 25056
rect 36580 24992 36596 25056
rect 36660 24992 36676 25056
rect 36740 24992 36756 25056
rect 36820 24992 36828 25056
rect 36508 23968 36828 24992
rect 36508 23904 36516 23968
rect 36580 23904 36596 23968
rect 36660 23904 36676 23968
rect 36740 23904 36756 23968
rect 36820 23904 36828 23968
rect 36508 22880 36828 23904
rect 36508 22816 36516 22880
rect 36580 22816 36596 22880
rect 36660 22816 36676 22880
rect 36740 22816 36756 22880
rect 36820 22816 36828 22880
rect 36508 21792 36828 22816
rect 36508 21728 36516 21792
rect 36580 21728 36596 21792
rect 36660 21728 36676 21792
rect 36740 21728 36756 21792
rect 36820 21728 36828 21792
rect 36508 20704 36828 21728
rect 36508 20640 36516 20704
rect 36580 20640 36596 20704
rect 36660 20640 36676 20704
rect 36740 20640 36756 20704
rect 36820 20640 36828 20704
rect 36508 19616 36828 20640
rect 36508 19552 36516 19616
rect 36580 19552 36596 19616
rect 36660 19552 36676 19616
rect 36740 19552 36756 19616
rect 36820 19552 36828 19616
rect 36508 18528 36828 19552
rect 36508 18464 36516 18528
rect 36580 18464 36596 18528
rect 36660 18464 36676 18528
rect 36740 18464 36756 18528
rect 36820 18464 36828 18528
rect 36508 17440 36828 18464
rect 36508 17376 36516 17440
rect 36580 17376 36596 17440
rect 36660 17376 36676 17440
rect 36740 17376 36756 17440
rect 36820 17376 36828 17440
rect 36508 16352 36828 17376
rect 36508 16288 36516 16352
rect 36580 16288 36596 16352
rect 36660 16288 36676 16352
rect 36740 16288 36756 16352
rect 36820 16288 36828 16352
rect 36508 15264 36828 16288
rect 36508 15200 36516 15264
rect 36580 15200 36596 15264
rect 36660 15200 36676 15264
rect 36740 15200 36756 15264
rect 36820 15200 36828 15264
rect 36508 14176 36828 15200
rect 36508 14112 36516 14176
rect 36580 14112 36596 14176
rect 36660 14112 36676 14176
rect 36740 14112 36756 14176
rect 36820 14112 36828 14176
rect 36508 13088 36828 14112
rect 36508 13024 36516 13088
rect 36580 13024 36596 13088
rect 36660 13024 36676 13088
rect 36740 13024 36756 13088
rect 36820 13024 36828 13088
rect 36508 12000 36828 13024
rect 36508 11936 36516 12000
rect 36580 11936 36596 12000
rect 36660 11936 36676 12000
rect 36740 11936 36756 12000
rect 36820 11936 36828 12000
rect 36508 10912 36828 11936
rect 36508 10848 36516 10912
rect 36580 10848 36596 10912
rect 36660 10848 36676 10912
rect 36740 10848 36756 10912
rect 36820 10848 36828 10912
rect 36508 9824 36828 10848
rect 36508 9760 36516 9824
rect 36580 9760 36596 9824
rect 36660 9760 36676 9824
rect 36740 9760 36756 9824
rect 36820 9760 36828 9824
rect 36508 8736 36828 9760
rect 36508 8672 36516 8736
rect 36580 8672 36596 8736
rect 36660 8672 36676 8736
rect 36740 8672 36756 8736
rect 36820 8672 36828 8736
rect 36508 7648 36828 8672
rect 36508 7584 36516 7648
rect 36580 7584 36596 7648
rect 36660 7584 36676 7648
rect 36740 7584 36756 7648
rect 36820 7584 36828 7648
rect 36508 6560 36828 7584
rect 36508 6496 36516 6560
rect 36580 6496 36596 6560
rect 36660 6496 36676 6560
rect 36740 6496 36756 6560
rect 36820 6496 36828 6560
rect 36508 6284 36828 6496
rect 36508 6048 36550 6284
rect 36786 6048 36828 6284
rect 36508 5472 36828 6048
rect 36508 5408 36516 5472
rect 36580 5408 36596 5472
rect 36660 5408 36676 5472
rect 36740 5408 36756 5472
rect 36820 5408 36828 5472
rect 36508 4384 36828 5408
rect 36508 4320 36516 4384
rect 36580 4320 36596 4384
rect 36660 4320 36676 4384
rect 36740 4320 36756 4384
rect 36820 4320 36828 4384
rect 36508 3296 36828 4320
rect 36508 3232 36516 3296
rect 36580 3232 36596 3296
rect 36660 3232 36676 3296
rect 36740 3232 36756 3296
rect 36820 3232 36828 3296
rect 36508 2208 36828 3232
rect 36508 2144 36516 2208
rect 36580 2144 36596 2208
rect 36660 2144 36676 2208
rect 36740 2144 36756 2208
rect 36820 2144 36828 2208
rect 36508 2128 36828 2144
rect 66568 77824 66888 77840
rect 66568 77760 66576 77824
rect 66640 77760 66656 77824
rect 66720 77760 66736 77824
rect 66800 77760 66816 77824
rect 66880 77760 66888 77824
rect 66568 76736 66888 77760
rect 66568 76672 66576 76736
rect 66640 76672 66656 76736
rect 66720 76672 66736 76736
rect 66800 76672 66816 76736
rect 66880 76672 66888 76736
rect 66568 75648 66888 76672
rect 66568 75584 66576 75648
rect 66640 75584 66656 75648
rect 66720 75584 66736 75648
rect 66800 75584 66816 75648
rect 66880 75584 66888 75648
rect 66568 74560 66888 75584
rect 66568 74496 66576 74560
rect 66640 74496 66656 74560
rect 66720 74496 66736 74560
rect 66800 74496 66816 74560
rect 66880 74496 66888 74560
rect 66568 73472 66888 74496
rect 66568 73408 66576 73472
rect 66640 73408 66656 73472
rect 66720 73408 66736 73472
rect 66800 73408 66816 73472
rect 66880 73408 66888 73472
rect 66568 72384 66888 73408
rect 66568 72320 66576 72384
rect 66640 72320 66656 72384
rect 66720 72320 66736 72384
rect 66800 72320 66816 72384
rect 66880 72320 66888 72384
rect 66568 71296 66888 72320
rect 66568 71232 66576 71296
rect 66640 71232 66656 71296
rect 66720 71232 66736 71296
rect 66800 71232 66816 71296
rect 66880 71232 66888 71296
rect 66568 70208 66888 71232
rect 66568 70144 66576 70208
rect 66640 70144 66656 70208
rect 66720 70144 66736 70208
rect 66800 70144 66816 70208
rect 66880 70144 66888 70208
rect 66568 69120 66888 70144
rect 66568 69056 66576 69120
rect 66640 69056 66656 69120
rect 66720 69056 66736 69120
rect 66800 69056 66816 69120
rect 66880 69056 66888 69120
rect 66568 68032 66888 69056
rect 66568 67968 66576 68032
rect 66640 67968 66656 68032
rect 66720 67968 66736 68032
rect 66800 67968 66816 68032
rect 66880 67968 66888 68032
rect 66568 66944 66888 67968
rect 66568 66880 66576 66944
rect 66640 66896 66656 66944
rect 66720 66896 66736 66944
rect 66800 66896 66816 66944
rect 66880 66880 66888 66944
rect 66568 66660 66610 66880
rect 66846 66660 66888 66880
rect 66568 65856 66888 66660
rect 66568 65792 66576 65856
rect 66640 65792 66656 65856
rect 66720 65792 66736 65856
rect 66800 65792 66816 65856
rect 66880 65792 66888 65856
rect 66568 64768 66888 65792
rect 66568 64704 66576 64768
rect 66640 64704 66656 64768
rect 66720 64704 66736 64768
rect 66800 64704 66816 64768
rect 66880 64704 66888 64768
rect 66568 63680 66888 64704
rect 66568 63616 66576 63680
rect 66640 63616 66656 63680
rect 66720 63616 66736 63680
rect 66800 63616 66816 63680
rect 66880 63616 66888 63680
rect 66568 62592 66888 63616
rect 66568 62528 66576 62592
rect 66640 62528 66656 62592
rect 66720 62528 66736 62592
rect 66800 62528 66816 62592
rect 66880 62528 66888 62592
rect 66568 61504 66888 62528
rect 66568 61440 66576 61504
rect 66640 61440 66656 61504
rect 66720 61440 66736 61504
rect 66800 61440 66816 61504
rect 66880 61440 66888 61504
rect 66568 60416 66888 61440
rect 66568 60352 66576 60416
rect 66640 60352 66656 60416
rect 66720 60352 66736 60416
rect 66800 60352 66816 60416
rect 66880 60352 66888 60416
rect 66568 59328 66888 60352
rect 66568 59264 66576 59328
rect 66640 59264 66656 59328
rect 66720 59264 66736 59328
rect 66800 59264 66816 59328
rect 66880 59264 66888 59328
rect 66568 58240 66888 59264
rect 66568 58176 66576 58240
rect 66640 58176 66656 58240
rect 66720 58176 66736 58240
rect 66800 58176 66816 58240
rect 66880 58176 66888 58240
rect 66568 57152 66888 58176
rect 66568 57088 66576 57152
rect 66640 57088 66656 57152
rect 66720 57088 66736 57152
rect 66800 57088 66816 57152
rect 66880 57088 66888 57152
rect 66568 56064 66888 57088
rect 66568 56000 66576 56064
rect 66640 56000 66656 56064
rect 66720 56000 66736 56064
rect 66800 56000 66816 56064
rect 66880 56000 66888 56064
rect 66568 54976 66888 56000
rect 66568 54912 66576 54976
rect 66640 54912 66656 54976
rect 66720 54912 66736 54976
rect 66800 54912 66816 54976
rect 66880 54912 66888 54976
rect 66568 53888 66888 54912
rect 66568 53824 66576 53888
rect 66640 53824 66656 53888
rect 66720 53824 66736 53888
rect 66800 53824 66816 53888
rect 66880 53824 66888 53888
rect 66568 52800 66888 53824
rect 66568 52736 66576 52800
rect 66640 52736 66656 52800
rect 66720 52736 66736 52800
rect 66800 52736 66816 52800
rect 66880 52736 66888 52800
rect 66568 51712 66888 52736
rect 66568 51648 66576 51712
rect 66640 51648 66656 51712
rect 66720 51648 66736 51712
rect 66800 51648 66816 51712
rect 66880 51648 66888 51712
rect 66568 50624 66888 51648
rect 66568 50560 66576 50624
rect 66640 50560 66656 50624
rect 66720 50560 66736 50624
rect 66800 50560 66816 50624
rect 66880 50560 66888 50624
rect 66568 49536 66888 50560
rect 66568 49472 66576 49536
rect 66640 49472 66656 49536
rect 66720 49472 66736 49536
rect 66800 49472 66816 49536
rect 66880 49472 66888 49536
rect 66568 48448 66888 49472
rect 66568 48384 66576 48448
rect 66640 48384 66656 48448
rect 66720 48384 66736 48448
rect 66800 48384 66816 48448
rect 66880 48384 66888 48448
rect 66568 47360 66888 48384
rect 66568 47296 66576 47360
rect 66640 47296 66656 47360
rect 66720 47296 66736 47360
rect 66800 47296 66816 47360
rect 66880 47296 66888 47360
rect 66568 46272 66888 47296
rect 66568 46208 66576 46272
rect 66640 46208 66656 46272
rect 66720 46208 66736 46272
rect 66800 46208 66816 46272
rect 66880 46208 66888 46272
rect 66568 45184 66888 46208
rect 66568 45120 66576 45184
rect 66640 45120 66656 45184
rect 66720 45120 66736 45184
rect 66800 45120 66816 45184
rect 66880 45120 66888 45184
rect 66568 44096 66888 45120
rect 66568 44032 66576 44096
rect 66640 44032 66656 44096
rect 66720 44032 66736 44096
rect 66800 44032 66816 44096
rect 66880 44032 66888 44096
rect 66568 43008 66888 44032
rect 66568 42944 66576 43008
rect 66640 42944 66656 43008
rect 66720 42944 66736 43008
rect 66800 42944 66816 43008
rect 66880 42944 66888 43008
rect 66568 41920 66888 42944
rect 66568 41856 66576 41920
rect 66640 41856 66656 41920
rect 66720 41856 66736 41920
rect 66800 41856 66816 41920
rect 66880 41856 66888 41920
rect 66568 40832 66888 41856
rect 66568 40768 66576 40832
rect 66640 40768 66656 40832
rect 66720 40768 66736 40832
rect 66800 40768 66816 40832
rect 66880 40768 66888 40832
rect 66568 39744 66888 40768
rect 66568 39680 66576 39744
rect 66640 39680 66656 39744
rect 66720 39680 66736 39744
rect 66800 39680 66816 39744
rect 66880 39680 66888 39744
rect 66568 38656 66888 39680
rect 66568 38592 66576 38656
rect 66640 38592 66656 38656
rect 66720 38592 66736 38656
rect 66800 38592 66816 38656
rect 66880 38592 66888 38656
rect 66568 37568 66888 38592
rect 66568 37504 66576 37568
rect 66640 37504 66656 37568
rect 66720 37504 66736 37568
rect 66800 37504 66816 37568
rect 66880 37504 66888 37568
rect 66568 36480 66888 37504
rect 66568 36416 66576 36480
rect 66640 36416 66656 36480
rect 66720 36416 66736 36480
rect 66800 36416 66816 36480
rect 66880 36416 66888 36480
rect 66568 36260 66888 36416
rect 66568 36024 66610 36260
rect 66846 36024 66888 36260
rect 66568 35392 66888 36024
rect 66568 35328 66576 35392
rect 66640 35328 66656 35392
rect 66720 35328 66736 35392
rect 66800 35328 66816 35392
rect 66880 35328 66888 35392
rect 66568 34304 66888 35328
rect 66568 34240 66576 34304
rect 66640 34240 66656 34304
rect 66720 34240 66736 34304
rect 66800 34240 66816 34304
rect 66880 34240 66888 34304
rect 66568 33216 66888 34240
rect 66568 33152 66576 33216
rect 66640 33152 66656 33216
rect 66720 33152 66736 33216
rect 66800 33152 66816 33216
rect 66880 33152 66888 33216
rect 66568 32128 66888 33152
rect 66568 32064 66576 32128
rect 66640 32064 66656 32128
rect 66720 32064 66736 32128
rect 66800 32064 66816 32128
rect 66880 32064 66888 32128
rect 66568 31040 66888 32064
rect 66568 30976 66576 31040
rect 66640 30976 66656 31040
rect 66720 30976 66736 31040
rect 66800 30976 66816 31040
rect 66880 30976 66888 31040
rect 66568 29952 66888 30976
rect 66568 29888 66576 29952
rect 66640 29888 66656 29952
rect 66720 29888 66736 29952
rect 66800 29888 66816 29952
rect 66880 29888 66888 29952
rect 66568 28864 66888 29888
rect 66568 28800 66576 28864
rect 66640 28800 66656 28864
rect 66720 28800 66736 28864
rect 66800 28800 66816 28864
rect 66880 28800 66888 28864
rect 66568 27776 66888 28800
rect 66568 27712 66576 27776
rect 66640 27712 66656 27776
rect 66720 27712 66736 27776
rect 66800 27712 66816 27776
rect 66880 27712 66888 27776
rect 66568 26688 66888 27712
rect 66568 26624 66576 26688
rect 66640 26624 66656 26688
rect 66720 26624 66736 26688
rect 66800 26624 66816 26688
rect 66880 26624 66888 26688
rect 66568 25600 66888 26624
rect 66568 25536 66576 25600
rect 66640 25536 66656 25600
rect 66720 25536 66736 25600
rect 66800 25536 66816 25600
rect 66880 25536 66888 25600
rect 66568 24512 66888 25536
rect 66568 24448 66576 24512
rect 66640 24448 66656 24512
rect 66720 24448 66736 24512
rect 66800 24448 66816 24512
rect 66880 24448 66888 24512
rect 66568 23424 66888 24448
rect 66568 23360 66576 23424
rect 66640 23360 66656 23424
rect 66720 23360 66736 23424
rect 66800 23360 66816 23424
rect 66880 23360 66888 23424
rect 66568 22336 66888 23360
rect 66568 22272 66576 22336
rect 66640 22272 66656 22336
rect 66720 22272 66736 22336
rect 66800 22272 66816 22336
rect 66880 22272 66888 22336
rect 66568 21248 66888 22272
rect 66568 21184 66576 21248
rect 66640 21184 66656 21248
rect 66720 21184 66736 21248
rect 66800 21184 66816 21248
rect 66880 21184 66888 21248
rect 66568 20160 66888 21184
rect 66568 20096 66576 20160
rect 66640 20096 66656 20160
rect 66720 20096 66736 20160
rect 66800 20096 66816 20160
rect 66880 20096 66888 20160
rect 66568 19072 66888 20096
rect 66568 19008 66576 19072
rect 66640 19008 66656 19072
rect 66720 19008 66736 19072
rect 66800 19008 66816 19072
rect 66880 19008 66888 19072
rect 66568 17984 66888 19008
rect 66568 17920 66576 17984
rect 66640 17920 66656 17984
rect 66720 17920 66736 17984
rect 66800 17920 66816 17984
rect 66880 17920 66888 17984
rect 66568 16896 66888 17920
rect 66568 16832 66576 16896
rect 66640 16832 66656 16896
rect 66720 16832 66736 16896
rect 66800 16832 66816 16896
rect 66880 16832 66888 16896
rect 66568 15808 66888 16832
rect 66568 15744 66576 15808
rect 66640 15744 66656 15808
rect 66720 15744 66736 15808
rect 66800 15744 66816 15808
rect 66880 15744 66888 15808
rect 66568 14720 66888 15744
rect 66568 14656 66576 14720
rect 66640 14656 66656 14720
rect 66720 14656 66736 14720
rect 66800 14656 66816 14720
rect 66880 14656 66888 14720
rect 66568 13632 66888 14656
rect 66568 13568 66576 13632
rect 66640 13568 66656 13632
rect 66720 13568 66736 13632
rect 66800 13568 66816 13632
rect 66880 13568 66888 13632
rect 66568 12544 66888 13568
rect 66568 12480 66576 12544
rect 66640 12480 66656 12544
rect 66720 12480 66736 12544
rect 66800 12480 66816 12544
rect 66880 12480 66888 12544
rect 66568 11456 66888 12480
rect 66568 11392 66576 11456
rect 66640 11392 66656 11456
rect 66720 11392 66736 11456
rect 66800 11392 66816 11456
rect 66880 11392 66888 11456
rect 66568 10368 66888 11392
rect 66568 10304 66576 10368
rect 66640 10304 66656 10368
rect 66720 10304 66736 10368
rect 66800 10304 66816 10368
rect 66880 10304 66888 10368
rect 66568 9280 66888 10304
rect 66568 9216 66576 9280
rect 66640 9216 66656 9280
rect 66720 9216 66736 9280
rect 66800 9216 66816 9280
rect 66880 9216 66888 9280
rect 66568 8192 66888 9216
rect 66568 8128 66576 8192
rect 66640 8128 66656 8192
rect 66720 8128 66736 8192
rect 66800 8128 66816 8192
rect 66880 8128 66888 8192
rect 66568 7104 66888 8128
rect 66568 7040 66576 7104
rect 66640 7040 66656 7104
rect 66720 7040 66736 7104
rect 66800 7040 66816 7104
rect 66880 7040 66888 7104
rect 66568 6016 66888 7040
rect 66568 5952 66576 6016
rect 66640 5952 66656 6016
rect 66720 5952 66736 6016
rect 66800 5952 66816 6016
rect 66880 5952 66888 6016
rect 66568 5624 66888 5952
rect 66568 5388 66610 5624
rect 66846 5388 66888 5624
rect 66568 4928 66888 5388
rect 66568 4864 66576 4928
rect 66640 4864 66656 4928
rect 66720 4864 66736 4928
rect 66800 4864 66816 4928
rect 66880 4864 66888 4928
rect 66568 3840 66888 4864
rect 66568 3776 66576 3840
rect 66640 3776 66656 3840
rect 66720 3776 66736 3840
rect 66800 3776 66816 3840
rect 66880 3776 66888 3840
rect 66568 2752 66888 3776
rect 66568 2688 66576 2752
rect 66640 2688 66656 2752
rect 66720 2688 66736 2752
rect 66800 2688 66816 2752
rect 66880 2688 66888 2752
rect 66568 2128 66888 2688
rect 67228 77280 67548 77840
rect 67228 77216 67236 77280
rect 67300 77216 67316 77280
rect 67380 77216 67396 77280
rect 67460 77216 67476 77280
rect 67540 77216 67548 77280
rect 67228 76192 67548 77216
rect 67228 76128 67236 76192
rect 67300 76128 67316 76192
rect 67380 76128 67396 76192
rect 67460 76128 67476 76192
rect 67540 76128 67548 76192
rect 67228 75104 67548 76128
rect 67228 75040 67236 75104
rect 67300 75040 67316 75104
rect 67380 75040 67396 75104
rect 67460 75040 67476 75104
rect 67540 75040 67548 75104
rect 67228 74016 67548 75040
rect 67228 73952 67236 74016
rect 67300 73952 67316 74016
rect 67380 73952 67396 74016
rect 67460 73952 67476 74016
rect 67540 73952 67548 74016
rect 67228 72928 67548 73952
rect 67228 72864 67236 72928
rect 67300 72864 67316 72928
rect 67380 72864 67396 72928
rect 67460 72864 67476 72928
rect 67540 72864 67548 72928
rect 67228 71840 67548 72864
rect 67228 71776 67236 71840
rect 67300 71776 67316 71840
rect 67380 71776 67396 71840
rect 67460 71776 67476 71840
rect 67540 71776 67548 71840
rect 67228 70752 67548 71776
rect 67228 70688 67236 70752
rect 67300 70688 67316 70752
rect 67380 70688 67396 70752
rect 67460 70688 67476 70752
rect 67540 70688 67548 70752
rect 67228 69664 67548 70688
rect 67228 69600 67236 69664
rect 67300 69600 67316 69664
rect 67380 69600 67396 69664
rect 67460 69600 67476 69664
rect 67540 69600 67548 69664
rect 67228 68576 67548 69600
rect 67228 68512 67236 68576
rect 67300 68512 67316 68576
rect 67380 68512 67396 68576
rect 67460 68512 67476 68576
rect 67540 68512 67548 68576
rect 67228 67556 67548 68512
rect 67228 67488 67270 67556
rect 67506 67488 67548 67556
rect 67228 67424 67236 67488
rect 67540 67424 67548 67488
rect 67228 67320 67270 67424
rect 67506 67320 67548 67424
rect 67228 66400 67548 67320
rect 67228 66336 67236 66400
rect 67300 66336 67316 66400
rect 67380 66336 67396 66400
rect 67460 66336 67476 66400
rect 67540 66336 67548 66400
rect 67228 65312 67548 66336
rect 67228 65248 67236 65312
rect 67300 65248 67316 65312
rect 67380 65248 67396 65312
rect 67460 65248 67476 65312
rect 67540 65248 67548 65312
rect 67228 64224 67548 65248
rect 67228 64160 67236 64224
rect 67300 64160 67316 64224
rect 67380 64160 67396 64224
rect 67460 64160 67476 64224
rect 67540 64160 67548 64224
rect 67228 63136 67548 64160
rect 67228 63072 67236 63136
rect 67300 63072 67316 63136
rect 67380 63072 67396 63136
rect 67460 63072 67476 63136
rect 67540 63072 67548 63136
rect 67228 62048 67548 63072
rect 67228 61984 67236 62048
rect 67300 61984 67316 62048
rect 67380 61984 67396 62048
rect 67460 61984 67476 62048
rect 67540 61984 67548 62048
rect 67228 60960 67548 61984
rect 67228 60896 67236 60960
rect 67300 60896 67316 60960
rect 67380 60896 67396 60960
rect 67460 60896 67476 60960
rect 67540 60896 67548 60960
rect 67228 59872 67548 60896
rect 67228 59808 67236 59872
rect 67300 59808 67316 59872
rect 67380 59808 67396 59872
rect 67460 59808 67476 59872
rect 67540 59808 67548 59872
rect 67228 58784 67548 59808
rect 67228 58720 67236 58784
rect 67300 58720 67316 58784
rect 67380 58720 67396 58784
rect 67460 58720 67476 58784
rect 67540 58720 67548 58784
rect 67228 57696 67548 58720
rect 67228 57632 67236 57696
rect 67300 57632 67316 57696
rect 67380 57632 67396 57696
rect 67460 57632 67476 57696
rect 67540 57632 67548 57696
rect 67228 56608 67548 57632
rect 67228 56544 67236 56608
rect 67300 56544 67316 56608
rect 67380 56544 67396 56608
rect 67460 56544 67476 56608
rect 67540 56544 67548 56608
rect 67228 55520 67548 56544
rect 67228 55456 67236 55520
rect 67300 55456 67316 55520
rect 67380 55456 67396 55520
rect 67460 55456 67476 55520
rect 67540 55456 67548 55520
rect 67228 54432 67548 55456
rect 67228 54368 67236 54432
rect 67300 54368 67316 54432
rect 67380 54368 67396 54432
rect 67460 54368 67476 54432
rect 67540 54368 67548 54432
rect 67228 53344 67548 54368
rect 67228 53280 67236 53344
rect 67300 53280 67316 53344
rect 67380 53280 67396 53344
rect 67460 53280 67476 53344
rect 67540 53280 67548 53344
rect 67228 52256 67548 53280
rect 67228 52192 67236 52256
rect 67300 52192 67316 52256
rect 67380 52192 67396 52256
rect 67460 52192 67476 52256
rect 67540 52192 67548 52256
rect 67228 51168 67548 52192
rect 67228 51104 67236 51168
rect 67300 51104 67316 51168
rect 67380 51104 67396 51168
rect 67460 51104 67476 51168
rect 67540 51104 67548 51168
rect 67228 50080 67548 51104
rect 67228 50016 67236 50080
rect 67300 50016 67316 50080
rect 67380 50016 67396 50080
rect 67460 50016 67476 50080
rect 67540 50016 67548 50080
rect 67228 48992 67548 50016
rect 67228 48928 67236 48992
rect 67300 48928 67316 48992
rect 67380 48928 67396 48992
rect 67460 48928 67476 48992
rect 67540 48928 67548 48992
rect 67228 47904 67548 48928
rect 67228 47840 67236 47904
rect 67300 47840 67316 47904
rect 67380 47840 67396 47904
rect 67460 47840 67476 47904
rect 67540 47840 67548 47904
rect 67228 46816 67548 47840
rect 67228 46752 67236 46816
rect 67300 46752 67316 46816
rect 67380 46752 67396 46816
rect 67460 46752 67476 46816
rect 67540 46752 67548 46816
rect 67228 45728 67548 46752
rect 67228 45664 67236 45728
rect 67300 45664 67316 45728
rect 67380 45664 67396 45728
rect 67460 45664 67476 45728
rect 67540 45664 67548 45728
rect 67228 44640 67548 45664
rect 67228 44576 67236 44640
rect 67300 44576 67316 44640
rect 67380 44576 67396 44640
rect 67460 44576 67476 44640
rect 67540 44576 67548 44640
rect 67228 43552 67548 44576
rect 67228 43488 67236 43552
rect 67300 43488 67316 43552
rect 67380 43488 67396 43552
rect 67460 43488 67476 43552
rect 67540 43488 67548 43552
rect 67228 42464 67548 43488
rect 67228 42400 67236 42464
rect 67300 42400 67316 42464
rect 67380 42400 67396 42464
rect 67460 42400 67476 42464
rect 67540 42400 67548 42464
rect 67228 41376 67548 42400
rect 67228 41312 67236 41376
rect 67300 41312 67316 41376
rect 67380 41312 67396 41376
rect 67460 41312 67476 41376
rect 67540 41312 67548 41376
rect 67228 40288 67548 41312
rect 67228 40224 67236 40288
rect 67300 40224 67316 40288
rect 67380 40224 67396 40288
rect 67460 40224 67476 40288
rect 67540 40224 67548 40288
rect 67228 39200 67548 40224
rect 67228 39136 67236 39200
rect 67300 39136 67316 39200
rect 67380 39136 67396 39200
rect 67460 39136 67476 39200
rect 67540 39136 67548 39200
rect 67228 38112 67548 39136
rect 67228 38048 67236 38112
rect 67300 38048 67316 38112
rect 67380 38048 67396 38112
rect 67460 38048 67476 38112
rect 67540 38048 67548 38112
rect 67228 37024 67548 38048
rect 67228 36960 67236 37024
rect 67300 36960 67316 37024
rect 67380 36960 67396 37024
rect 67460 36960 67476 37024
rect 67540 36960 67548 37024
rect 67228 36920 67548 36960
rect 67228 36684 67270 36920
rect 67506 36684 67548 36920
rect 67228 35936 67548 36684
rect 67228 35872 67236 35936
rect 67300 35872 67316 35936
rect 67380 35872 67396 35936
rect 67460 35872 67476 35936
rect 67540 35872 67548 35936
rect 67228 34848 67548 35872
rect 67228 34784 67236 34848
rect 67300 34784 67316 34848
rect 67380 34784 67396 34848
rect 67460 34784 67476 34848
rect 67540 34784 67548 34848
rect 67228 33760 67548 34784
rect 67228 33696 67236 33760
rect 67300 33696 67316 33760
rect 67380 33696 67396 33760
rect 67460 33696 67476 33760
rect 67540 33696 67548 33760
rect 67228 32672 67548 33696
rect 67228 32608 67236 32672
rect 67300 32608 67316 32672
rect 67380 32608 67396 32672
rect 67460 32608 67476 32672
rect 67540 32608 67548 32672
rect 67228 31584 67548 32608
rect 67228 31520 67236 31584
rect 67300 31520 67316 31584
rect 67380 31520 67396 31584
rect 67460 31520 67476 31584
rect 67540 31520 67548 31584
rect 67228 30496 67548 31520
rect 67228 30432 67236 30496
rect 67300 30432 67316 30496
rect 67380 30432 67396 30496
rect 67460 30432 67476 30496
rect 67540 30432 67548 30496
rect 67228 29408 67548 30432
rect 67228 29344 67236 29408
rect 67300 29344 67316 29408
rect 67380 29344 67396 29408
rect 67460 29344 67476 29408
rect 67540 29344 67548 29408
rect 67228 28320 67548 29344
rect 67228 28256 67236 28320
rect 67300 28256 67316 28320
rect 67380 28256 67396 28320
rect 67460 28256 67476 28320
rect 67540 28256 67548 28320
rect 67228 27232 67548 28256
rect 67228 27168 67236 27232
rect 67300 27168 67316 27232
rect 67380 27168 67396 27232
rect 67460 27168 67476 27232
rect 67540 27168 67548 27232
rect 67228 26144 67548 27168
rect 67228 26080 67236 26144
rect 67300 26080 67316 26144
rect 67380 26080 67396 26144
rect 67460 26080 67476 26144
rect 67540 26080 67548 26144
rect 67228 25056 67548 26080
rect 67228 24992 67236 25056
rect 67300 24992 67316 25056
rect 67380 24992 67396 25056
rect 67460 24992 67476 25056
rect 67540 24992 67548 25056
rect 67228 23968 67548 24992
rect 67228 23904 67236 23968
rect 67300 23904 67316 23968
rect 67380 23904 67396 23968
rect 67460 23904 67476 23968
rect 67540 23904 67548 23968
rect 67228 22880 67548 23904
rect 67228 22816 67236 22880
rect 67300 22816 67316 22880
rect 67380 22816 67396 22880
rect 67460 22816 67476 22880
rect 67540 22816 67548 22880
rect 67228 21792 67548 22816
rect 67228 21728 67236 21792
rect 67300 21728 67316 21792
rect 67380 21728 67396 21792
rect 67460 21728 67476 21792
rect 67540 21728 67548 21792
rect 67228 20704 67548 21728
rect 67228 20640 67236 20704
rect 67300 20640 67316 20704
rect 67380 20640 67396 20704
rect 67460 20640 67476 20704
rect 67540 20640 67548 20704
rect 67228 19616 67548 20640
rect 67228 19552 67236 19616
rect 67300 19552 67316 19616
rect 67380 19552 67396 19616
rect 67460 19552 67476 19616
rect 67540 19552 67548 19616
rect 67228 18528 67548 19552
rect 67228 18464 67236 18528
rect 67300 18464 67316 18528
rect 67380 18464 67396 18528
rect 67460 18464 67476 18528
rect 67540 18464 67548 18528
rect 67228 17440 67548 18464
rect 67228 17376 67236 17440
rect 67300 17376 67316 17440
rect 67380 17376 67396 17440
rect 67460 17376 67476 17440
rect 67540 17376 67548 17440
rect 67228 16352 67548 17376
rect 67228 16288 67236 16352
rect 67300 16288 67316 16352
rect 67380 16288 67396 16352
rect 67460 16288 67476 16352
rect 67540 16288 67548 16352
rect 67228 15264 67548 16288
rect 67228 15200 67236 15264
rect 67300 15200 67316 15264
rect 67380 15200 67396 15264
rect 67460 15200 67476 15264
rect 67540 15200 67548 15264
rect 67228 14176 67548 15200
rect 67228 14112 67236 14176
rect 67300 14112 67316 14176
rect 67380 14112 67396 14176
rect 67460 14112 67476 14176
rect 67540 14112 67548 14176
rect 67228 13088 67548 14112
rect 67228 13024 67236 13088
rect 67300 13024 67316 13088
rect 67380 13024 67396 13088
rect 67460 13024 67476 13088
rect 67540 13024 67548 13088
rect 67228 12000 67548 13024
rect 67228 11936 67236 12000
rect 67300 11936 67316 12000
rect 67380 11936 67396 12000
rect 67460 11936 67476 12000
rect 67540 11936 67548 12000
rect 67228 10912 67548 11936
rect 67228 10848 67236 10912
rect 67300 10848 67316 10912
rect 67380 10848 67396 10912
rect 67460 10848 67476 10912
rect 67540 10848 67548 10912
rect 67228 9824 67548 10848
rect 67228 9760 67236 9824
rect 67300 9760 67316 9824
rect 67380 9760 67396 9824
rect 67460 9760 67476 9824
rect 67540 9760 67548 9824
rect 67228 8736 67548 9760
rect 67228 8672 67236 8736
rect 67300 8672 67316 8736
rect 67380 8672 67396 8736
rect 67460 8672 67476 8736
rect 67540 8672 67548 8736
rect 67228 7648 67548 8672
rect 67228 7584 67236 7648
rect 67300 7584 67316 7648
rect 67380 7584 67396 7648
rect 67460 7584 67476 7648
rect 67540 7584 67548 7648
rect 67228 6560 67548 7584
rect 67228 6496 67236 6560
rect 67300 6496 67316 6560
rect 67380 6496 67396 6560
rect 67460 6496 67476 6560
rect 67540 6496 67548 6560
rect 67228 6284 67548 6496
rect 67228 6048 67270 6284
rect 67506 6048 67548 6284
rect 67228 5472 67548 6048
rect 67228 5408 67236 5472
rect 67300 5408 67316 5472
rect 67380 5408 67396 5472
rect 67460 5408 67476 5472
rect 67540 5408 67548 5472
rect 67228 4384 67548 5408
rect 67228 4320 67236 4384
rect 67300 4320 67316 4384
rect 67380 4320 67396 4384
rect 67460 4320 67476 4384
rect 67540 4320 67548 4384
rect 67228 3296 67548 4320
rect 67228 3232 67236 3296
rect 67300 3232 67316 3296
rect 67380 3232 67396 3296
rect 67460 3232 67476 3296
rect 67540 3232 67548 3296
rect 67228 2208 67548 3232
rect 67228 2144 67236 2208
rect 67300 2144 67316 2208
rect 67380 2144 67396 2208
rect 67460 2144 67476 2208
rect 67540 2144 67548 2208
rect 67228 2128 67548 2144
<< via4 >>
rect 5170 66880 5200 66896
rect 5200 66880 5216 66896
rect 5216 66880 5280 66896
rect 5280 66880 5296 66896
rect 5296 66880 5360 66896
rect 5360 66880 5376 66896
rect 5376 66880 5406 66896
rect 5170 66660 5406 66880
rect 5170 36024 5406 36260
rect 5170 5388 5406 5624
rect 5830 67488 6066 67556
rect 5830 67424 5860 67488
rect 5860 67424 5876 67488
rect 5876 67424 5940 67488
rect 5940 67424 5956 67488
rect 5956 67424 6020 67488
rect 6020 67424 6036 67488
rect 6036 67424 6066 67488
rect 5830 67320 6066 67424
rect 5830 36684 6066 36920
rect 5830 6048 6066 6284
rect 35890 66880 35920 66896
rect 35920 66880 35936 66896
rect 35936 66880 36000 66896
rect 36000 66880 36016 66896
rect 36016 66880 36080 66896
rect 36080 66880 36096 66896
rect 36096 66880 36126 66896
rect 35890 66660 36126 66880
rect 35890 36024 36126 36260
rect 35890 5388 36126 5624
rect 36550 67488 36786 67556
rect 36550 67424 36580 67488
rect 36580 67424 36596 67488
rect 36596 67424 36660 67488
rect 36660 67424 36676 67488
rect 36676 67424 36740 67488
rect 36740 67424 36756 67488
rect 36756 67424 36786 67488
rect 36550 67320 36786 67424
rect 36550 36684 36786 36920
rect 36550 6048 36786 6284
rect 66610 66880 66640 66896
rect 66640 66880 66656 66896
rect 66656 66880 66720 66896
rect 66720 66880 66736 66896
rect 66736 66880 66800 66896
rect 66800 66880 66816 66896
rect 66816 66880 66846 66896
rect 66610 66660 66846 66880
rect 66610 36024 66846 36260
rect 66610 5388 66846 5624
rect 67270 67488 67506 67556
rect 67270 67424 67300 67488
rect 67300 67424 67316 67488
rect 67316 67424 67380 67488
rect 67380 67424 67396 67488
rect 67396 67424 67460 67488
rect 67460 67424 67476 67488
rect 67476 67424 67506 67488
rect 67270 67320 67506 67424
rect 67270 36684 67506 36920
rect 67270 6048 67506 6284
<< metal5 >>
rect 1976 67556 77972 67598
rect 1976 67320 5830 67556
rect 6066 67320 36550 67556
rect 36786 67320 67270 67556
rect 67506 67320 77972 67556
rect 1976 67278 77972 67320
rect 1976 66896 77972 66938
rect 1976 66660 5170 66896
rect 5406 66660 35890 66896
rect 36126 66660 66610 66896
rect 66846 66660 77972 66896
rect 1976 66618 77972 66660
rect 1976 36920 77972 36962
rect 1976 36684 5830 36920
rect 6066 36684 36550 36920
rect 36786 36684 67270 36920
rect 67506 36684 77972 36920
rect 1976 36642 77972 36684
rect 1976 36260 77972 36302
rect 1976 36024 5170 36260
rect 5406 36024 35890 36260
rect 36126 36024 66610 36260
rect 66846 36024 77972 36260
rect 1976 35982 77972 36024
rect 1976 6284 77972 6326
rect 1976 6048 5830 6284
rect 6066 6048 36550 6284
rect 36786 6048 67270 6284
rect 67506 6048 77972 6284
rect 1976 6006 77972 6048
rect 1976 5624 77972 5666
rect 1976 5388 5170 5624
rect 5406 5388 35890 5624
rect 36126 5388 66610 5624
rect 66846 5388 77972 5624
rect 1976 5346 77972 5388
use sky130_fd_sc_hd__inv_2  _030_
timestamp 1
transform 1 0 74612 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _031_
timestamp 1
transform -1 0 58236 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _032_
timestamp 1
transform -1 0 59064 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _033_
timestamp 1
transform -1 0 75992 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _034_
timestamp 1
transform -1 0 75440 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _035_
timestamp 1
transform -1 0 72036 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _036_
timestamp 1
transform -1 0 76268 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _037_
timestamp 1
transform 1 0 57500 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _038_
timestamp 1
transform -1 0 58052 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _039_
timestamp 1
transform -1 0 57500 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _040_
timestamp 1
transform -1 0 56948 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _041_
timestamp 1
transform 1 0 59984 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _042_
timestamp 1
transform -1 0 60536 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _043_
timestamp 1
transform -1 0 61088 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _044_
timestamp 1
transform 1 0 64584 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _045_
timestamp 1
transform 1 0 60628 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _046_
timestamp 1
transform 1 0 64768 0 1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _047_
timestamp 1
transform -1 0 66240 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _048_
timestamp 1
transform -1 0 66332 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _049_
timestamp 1
transform 1 0 66240 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _050_
timestamp 1
transform 1 0 66516 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _051_
timestamp 1
transform -1 0 66792 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _052_
timestamp 1
transform 1 0 65412 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _053_
timestamp 1
transform 1 0 65688 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _054_
timestamp 1
transform -1 0 71484 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _055_
timestamp 1
transform 1 0 70564 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _056_
timestamp 1
transform -1 0 70932 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _057_
timestamp 1
transform -1 0 71944 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _058_
timestamp 1
transform 1 0 72588 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _059_
timestamp 1
transform -1 0 71484 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _060_
timestamp 1
transform -1 0 71576 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _061_
timestamp 1
transform -1 0 71208 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _062_
timestamp 1
transform 1 0 74244 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _064_
timestamp 1
transform -1 0 58420 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1
transform -1 0 62468 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _066_
timestamp 1
transform 1 0 61732 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _067_
timestamp 1
transform -1 0 67252 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _068_
timestamp 1
transform -1 0 67344 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _069_
timestamp 1
transform -1 0 66240 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1
transform 1 0 66792 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _071_
timestamp 1
transform -1 0 71116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _072_
timestamp 1
transform -1 0 76268 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 1
transform -1 0 71392 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 1
transform -1 0 76452 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _075_
timestamp 1
transform 1 0 57592 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _076_
timestamp 1
transform 1 0 56764 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _077_
timestamp 1
transform 1 0 56304 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _078_
timestamp 1
transform 1 0 60352 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _079_
timestamp 1
transform 1 0 61364 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _080_
timestamp 1
transform 1 0 65136 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _081_
timestamp 1
transform -1 0 68356 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _082_
timestamp 1
transform 1 0 64308 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _083_
timestamp 1
transform -1 0 68356 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _084_
timestamp 1
transform -1 0 71668 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _085_
timestamp 1
transform 1 0 74060 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _086_
timestamp 1
transform 1 0 70196 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _087_
timestamp 1
transform 1 0 74336 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1
transform -1 0 76360 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1
transform -1 0 76544 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform 1 0 65412 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1
transform -1 0 64768 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1
transform 1 0 67804 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 1
transform 1 0 67804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout6
timestamp 1
transform -1 0 72220 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 3404 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 4692 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 5796 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 7268 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 8372 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636968456
transform 1 0 9844 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636968456
transform 1 0 10948 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 12420 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636968456
transform 1 0 13524 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14996 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 16100 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 17572 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636968456
transform 1 0 18676 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636968456
transform 1 0 20148 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636968456
transform 1 0 21252 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_228
timestamp 1
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_234
timestamp 1636968456
transform 1 0 23552 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1
transform 1 0 24656 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636968456
transform 1 0 25300 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636968456
transform 1 0 26404 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636968456
transform 1 0 27876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636968456
transform 1 0 28980 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636968456
transform 1 0 30452 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636968456
transform 1 0 31556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 1
transform 1 0 33028 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_346
timestamp 1636968456
transform 1 0 33856 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_358
timestamp 1
transform 1 0 34960 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636968456
transform 1 0 35604 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636968456
transform 1 0 36708 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1
transform 1 0 37812 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1636968456
transform 1 0 38180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1636968456
transform 1 0 39284 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1
transform 1 0 40388 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1636968456
transform 1 0 40756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_433
timestamp 1
transform 1 0 41860 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_437
timestamp 1
transform 1 0 42228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1636968456
transform 1 0 43332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_461
timestamp 1
transform 1 0 44436 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_465
timestamp 1
transform 1 0 44804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1
transform 1 0 45540 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1636968456
transform 1 0 45908 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1636968456
transform 1 0 47012 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1
transform 1 0 48116 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1636968456
transform 1 0 48484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_517
timestamp 1636968456
transform 1 0 49588 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1
transform 1 0 50692 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_533
timestamp 1636968456
transform 1 0 51060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_545
timestamp 1
transform 1 0 52164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_549
timestamp 1
transform 1 0 52532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1
transform 1 0 53268 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_561
timestamp 1636968456
transform 1 0 53636 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_573
timestamp 1636968456
transform 1 0 54740 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1
transform 1 0 55844 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_589
timestamp 1636968456
transform 1 0 56212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_601
timestamp 1
transform 1 0 57316 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_612
timestamp 1
transform 1 0 58328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_617
timestamp 1
transform 1 0 58788 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_626
timestamp 1636968456
transform 1 0 59616 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_638
timestamp 1
transform 1 0 60720 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1636968456
transform 1 0 61364 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1636968456
transform 1 0 62468 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1
transform 1 0 63572 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1636968456
transform 1 0 63940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1636968456
transform 1 0 65044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1
transform 1 0 66148 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1636968456
transform 1 0 66516 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1636968456
transform 1 0 67620 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1
transform 1 0 68724 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_729
timestamp 1636968456
transform 1 0 69092 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_741
timestamp 1636968456
transform 1 0 70196 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1
transform 1 0 71300 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_757
timestamp 1636968456
transform 1 0 71668 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_769
timestamp 1636968456
transform 1 0 72772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 1
transform 1 0 73876 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_785
timestamp 1636968456
transform 1 0 74244 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_797
timestamp 1636968456
transform 1 0 75348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 1
transform 1 0 76452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_813
timestamp 1
transform 1 0 76820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_821
timestamp 1
transform 1 0 77556 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 2300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 3404 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 4508 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 5612 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 7084 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636968456
transform 1 0 7268 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 8372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636968456
transform 1 0 9476 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636968456
transform 1 0 10580 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1
transform 1 0 11684 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636968456
transform 1 0 12420 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636968456
transform 1 0 13524 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636968456
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636968456
transform 1 0 15732 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1
transform 1 0 16836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636968456
transform 1 0 17572 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636968456
transform 1 0 18676 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636968456
transform 1 0 19780 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636968456
transform 1 0 20884 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1
transform 1 0 21988 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636968456
transform 1 0 22724 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636968456
transform 1 0 23828 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636968456
transform 1 0 24932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636968456
transform 1 0 26036 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1
transform 1 0 27140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1
transform 1 0 27692 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636968456
transform 1 0 27876 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636968456
transform 1 0 28980 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636968456
transform 1 0 30084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636968456
transform 1 0 31188 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1
transform 1 0 32292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1
transform 1 0 32844 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636968456
transform 1 0 33028 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636968456
transform 1 0 34132 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636968456
transform 1 0 35236 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636968456
transform 1 0 36340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1
transform 1 0 37444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1
transform 1 0 37996 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636968456
transform 1 0 38180 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636968456
transform 1 0 39284 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636968456
transform 1 0 40388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636968456
transform 1 0 41492 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1
transform 1 0 42596 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1
transform 1 0 43148 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636968456
transform 1 0 43332 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636968456
transform 1 0 44436 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636968456
transform 1 0 45540 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636968456
transform 1 0 46644 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1
transform 1 0 47748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1
transform 1 0 48300 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636968456
transform 1 0 48484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636968456
transform 1 0 49588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636968456
transform 1 0 50692 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636968456
transform 1 0 51796 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1
transform 1 0 52900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1
transform 1 0 53452 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636968456
transform 1 0 53636 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636968456
transform 1 0 54740 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636968456
transform 1 0 55844 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636968456
transform 1 0 56948 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1
transform 1 0 58052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1
transform 1 0 58604 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636968456
transform 1 0 58788 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636968456
transform 1 0 59892 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636968456
transform 1 0 60996 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636968456
transform 1 0 62100 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 1
transform 1 0 63204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1
transform 1 0 63756 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636968456
transform 1 0 63940 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636968456
transform 1 0 65044 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636968456
transform 1 0 66148 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636968456
transform 1 0 67252 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1
transform 1 0 68356 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1
transform 1 0 68908 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636968456
transform 1 0 69092 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636968456
transform 1 0 70196 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636968456
transform 1 0 71300 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636968456
transform 1 0 72404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 1
transform 1 0 73508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 1
transform 1 0 74060 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636968456
transform 1 0 74244 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636968456
transform 1 0 75348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636968456
transform 1 0 76452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_821
timestamp 1
transform 1 0 77556 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 2300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 3404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 4692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636968456
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636968456
transform 1 0 6900 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636968456
transform 1 0 8004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1
transform 1 0 9108 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 9660 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636968456
transform 1 0 9844 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636968456
transform 1 0 10948 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636968456
transform 1 0 12052 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636968456
transform 1 0 13156 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1
transform 1 0 14260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 14812 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636968456
transform 1 0 14996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636968456
transform 1 0 16100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636968456
transform 1 0 17204 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636968456
transform 1 0 18308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1
transform 1 0 19412 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 19964 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636968456
transform 1 0 20148 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636968456
transform 1 0 21252 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636968456
transform 1 0 22356 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636968456
transform 1 0 23460 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1
transform 1 0 24564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 25116 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636968456
transform 1 0 25300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636968456
transform 1 0 26404 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636968456
transform 1 0 27508 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636968456
transform 1 0 28612 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1
transform 1 0 29716 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1
transform 1 0 30268 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636968456
transform 1 0 30452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636968456
transform 1 0 31556 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636968456
transform 1 0 32660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636968456
transform 1 0 33764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1
transform 1 0 34868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1
transform 1 0 35420 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636968456
transform 1 0 35604 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636968456
transform 1 0 36708 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636968456
transform 1 0 37812 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636968456
transform 1 0 38916 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1
transform 1 0 40020 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1
transform 1 0 40572 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636968456
transform 1 0 40756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636968456
transform 1 0 41860 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636968456
transform 1 0 42964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636968456
transform 1 0 44068 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1
transform 1 0 45172 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1
transform 1 0 45724 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636968456
transform 1 0 45908 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636968456
transform 1 0 47012 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636968456
transform 1 0 48116 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636968456
transform 1 0 49220 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1
transform 1 0 50324 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1
transform 1 0 50876 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636968456
transform 1 0 51060 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636968456
transform 1 0 52164 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636968456
transform 1 0 53268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636968456
transform 1 0 54372 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1
transform 1 0 55476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1
transform 1 0 56028 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636968456
transform 1 0 56212 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636968456
transform 1 0 57316 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636968456
transform 1 0 58420 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636968456
transform 1 0 59524 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1
transform 1 0 60628 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1
transform 1 0 61180 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636968456
transform 1 0 61364 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636968456
transform 1 0 62468 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636968456
transform 1 0 63572 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636968456
transform 1 0 64676 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1
transform 1 0 65780 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1
transform 1 0 66332 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636968456
transform 1 0 66516 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636968456
transform 1 0 67620 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636968456
transform 1 0 68724 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636968456
transform 1 0 69828 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1
transform 1 0 70932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1
transform 1 0 71484 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636968456
transform 1 0 71668 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636968456
transform 1 0 72772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636968456
transform 1 0 73876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636968456
transform 1 0 74980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1
transform 1 0 76084 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1
transform 1 0 76636 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_813
timestamp 1
transform 1 0 76820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_821
timestamp 1
transform 1 0 77556 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 2300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 3404 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 4508 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 5612 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1
transform 1 0 6716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636968456
transform 1 0 7268 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636968456
transform 1 0 8372 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636968456
transform 1 0 9476 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636968456
transform 1 0 10580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1
transform 1 0 11684 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636968456
transform 1 0 12420 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636968456
transform 1 0 13524 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636968456
transform 1 0 14628 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636968456
transform 1 0 15732 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1
transform 1 0 16836 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636968456
transform 1 0 17572 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636968456
transform 1 0 18676 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636968456
transform 1 0 19780 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636968456
transform 1 0 20884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1
transform 1 0 21988 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 22540 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636968456
transform 1 0 22724 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636968456
transform 1 0 23828 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636968456
transform 1 0 24932 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636968456
transform 1 0 26036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1
transform 1 0 27140 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1
transform 1 0 27692 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636968456
transform 1 0 27876 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636968456
transform 1 0 28980 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636968456
transform 1 0 30084 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636968456
transform 1 0 31188 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1
transform 1 0 32292 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1
transform 1 0 32844 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636968456
transform 1 0 33028 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636968456
transform 1 0 34132 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636968456
transform 1 0 35236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636968456
transform 1 0 36340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1
transform 1 0 37444 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1
transform 1 0 37996 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636968456
transform 1 0 38180 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636968456
transform 1 0 39284 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636968456
transform 1 0 40388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636968456
transform 1 0 41492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1
transform 1 0 42596 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1
transform 1 0 43148 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636968456
transform 1 0 43332 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636968456
transform 1 0 44436 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636968456
transform 1 0 45540 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636968456
transform 1 0 46644 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1
transform 1 0 47748 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1
transform 1 0 48300 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636968456
transform 1 0 48484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636968456
transform 1 0 49588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636968456
transform 1 0 50692 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636968456
transform 1 0 51796 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1
transform 1 0 52900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1
transform 1 0 53452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636968456
transform 1 0 53636 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636968456
transform 1 0 54740 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636968456
transform 1 0 55844 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636968456
transform 1 0 56948 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1
transform 1 0 58052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1
transform 1 0 58604 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636968456
transform 1 0 58788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636968456
transform 1 0 59892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636968456
transform 1 0 60996 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636968456
transform 1 0 62100 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1
transform 1 0 63204 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1
transform 1 0 63756 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636968456
transform 1 0 63940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636968456
transform 1 0 65044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636968456
transform 1 0 66148 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636968456
transform 1 0 67252 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1
transform 1 0 68356 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1
transform 1 0 68908 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636968456
transform 1 0 69092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636968456
transform 1 0 70196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636968456
transform 1 0 71300 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636968456
transform 1 0 72404 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1
transform 1 0 73508 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1
transform 1 0 74060 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636968456
transform 1 0 74244 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636968456
transform 1 0 75348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636968456
transform 1 0 76452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_821
timestamp 1
transform 1 0 77556 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 3404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 4692 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636968456
transform 1 0 5796 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636968456
transform 1 0 6900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636968456
transform 1 0 8004 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1
transform 1 0 9108 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 9660 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636968456
transform 1 0 9844 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636968456
transform 1 0 10948 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636968456
transform 1 0 12052 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636968456
transform 1 0 13156 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1
transform 1 0 14260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 14812 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14996 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636968456
transform 1 0 16100 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636968456
transform 1 0 17204 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636968456
transform 1 0 18308 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1
transform 1 0 19412 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 19964 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636968456
transform 1 0 20148 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636968456
transform 1 0 21252 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636968456
transform 1 0 22356 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636968456
transform 1 0 23460 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1
transform 1 0 24564 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 25116 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636968456
transform 1 0 25300 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636968456
transform 1 0 26404 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636968456
transform 1 0 27508 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636968456
transform 1 0 28612 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1
transform 1 0 29716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1
transform 1 0 30268 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636968456
transform 1 0 30452 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636968456
transform 1 0 31556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636968456
transform 1 0 32660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636968456
transform 1 0 33764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1
transform 1 0 34868 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1
transform 1 0 35420 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636968456
transform 1 0 35604 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636968456
transform 1 0 36708 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636968456
transform 1 0 37812 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636968456
transform 1 0 38916 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1
transform 1 0 40020 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1
transform 1 0 40572 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636968456
transform 1 0 40756 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636968456
transform 1 0 41860 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1636968456
transform 1 0 42964 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1636968456
transform 1 0 44068 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1
transform 1 0 45172 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1
transform 1 0 45724 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636968456
transform 1 0 45908 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636968456
transform 1 0 47012 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1636968456
transform 1 0 48116 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1636968456
transform 1 0 49220 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1
transform 1 0 50324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1
transform 1 0 50876 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636968456
transform 1 0 51060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636968456
transform 1 0 52164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1636968456
transform 1 0 53268 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1636968456
transform 1 0 54372 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1
transform 1 0 55476 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1
transform 1 0 56028 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636968456
transform 1 0 56212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636968456
transform 1 0 57316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1636968456
transform 1 0 58420 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1636968456
transform 1 0 59524 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1
transform 1 0 60628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1
transform 1 0 61180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636968456
transform 1 0 61364 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636968456
transform 1 0 62468 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1636968456
transform 1 0 63572 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1636968456
transform 1 0 64676 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1
transform 1 0 65780 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1
transform 1 0 66332 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636968456
transform 1 0 66516 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636968456
transform 1 0 67620 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1636968456
transform 1 0 68724 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1636968456
transform 1 0 69828 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1
transform 1 0 70932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1
transform 1 0 71484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636968456
transform 1 0 71668 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636968456
transform 1 0 72772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1636968456
transform 1 0 73876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1636968456
transform 1 0 74980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1
transform 1 0 76084 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1
transform 1 0 76636 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_813
timestamp 1
transform 1 0 76820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_821
timestamp 1
transform 1 0 77556 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636968456
transform 1 0 2300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636968456
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636968456
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636968456
transform 1 0 5612 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1
transform 1 0 6716 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 7084 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636968456
transform 1 0 7268 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636968456
transform 1 0 8372 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636968456
transform 1 0 9476 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636968456
transform 1 0 10580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1
transform 1 0 11684 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 12236 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636968456
transform 1 0 12420 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636968456
transform 1 0 13524 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636968456
transform 1 0 14628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636968456
transform 1 0 15732 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1
transform 1 0 16836 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636968456
transform 1 0 17572 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636968456
transform 1 0 18676 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636968456
transform 1 0 19780 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636968456
transform 1 0 20884 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1
transform 1 0 21988 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 22540 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636968456
transform 1 0 22724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636968456
transform 1 0 23828 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636968456
transform 1 0 24932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636968456
transform 1 0 26036 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1
transform 1 0 27140 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 27692 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636968456
transform 1 0 27876 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636968456
transform 1 0 28980 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636968456
transform 1 0 30084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636968456
transform 1 0 31188 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1
transform 1 0 32292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1
transform 1 0 32844 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636968456
transform 1 0 33028 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636968456
transform 1 0 34132 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636968456
transform 1 0 35236 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636968456
transform 1 0 36340 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1
transform 1 0 37444 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1
transform 1 0 37996 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636968456
transform 1 0 38180 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636968456
transform 1 0 39284 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636968456
transform 1 0 40388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636968456
transform 1 0 41492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1
transform 1 0 42596 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1
transform 1 0 43148 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1636968456
transform 1 0 43332 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1636968456
transform 1 0 44436 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1636968456
transform 1 0 45540 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1636968456
transform 1 0 46644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1
transform 1 0 47748 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1
transform 1 0 48300 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1636968456
transform 1 0 48484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1636968456
transform 1 0 49588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1636968456
transform 1 0 50692 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1636968456
transform 1 0 51796 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1
transform 1 0 52900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1
transform 1 0 53452 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1636968456
transform 1 0 53636 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1636968456
transform 1 0 54740 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1636968456
transform 1 0 55844 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1636968456
transform 1 0 56948 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1
transform 1 0 58052 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1
transform 1 0 58604 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1636968456
transform 1 0 58788 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1636968456
transform 1 0 59892 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1636968456
transform 1 0 60996 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1636968456
transform 1 0 62100 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1
transform 1 0 63204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1
transform 1 0 63756 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1636968456
transform 1 0 63940 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1636968456
transform 1 0 65044 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1636968456
transform 1 0 66148 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1636968456
transform 1 0 67252 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1
transform 1 0 68356 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1
transform 1 0 68908 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1636968456
transform 1 0 69092 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1636968456
transform 1 0 70196 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1636968456
transform 1 0 71300 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1636968456
transform 1 0 72404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1
transform 1 0 73508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1
transform 1 0 74060 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1636968456
transform 1 0 74244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1636968456
transform 1 0 75348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1636968456
transform 1 0 76452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_821
timestamp 1
transform 1 0 77556 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636968456
transform 1 0 2300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636968456
transform 1 0 3404 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 4508 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 4692 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636968456
transform 1 0 5796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636968456
transform 1 0 6900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636968456
transform 1 0 8004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1
transform 1 0 9108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636968456
transform 1 0 9844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636968456
transform 1 0 10948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636968456
transform 1 0 12052 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636968456
transform 1 0 13156 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1
transform 1 0 14260 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 14812 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636968456
transform 1 0 14996 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636968456
transform 1 0 16100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636968456
transform 1 0 17204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636968456
transform 1 0 18308 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1
transform 1 0 19412 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19964 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636968456
transform 1 0 20148 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636968456
transform 1 0 21252 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636968456
transform 1 0 22356 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636968456
transform 1 0 23460 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1
transform 1 0 24564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 25116 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636968456
transform 1 0 25300 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636968456
transform 1 0 26404 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636968456
transform 1 0 27508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636968456
transform 1 0 28612 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1
transform 1 0 29716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1
transform 1 0 30268 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636968456
transform 1 0 30452 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636968456
transform 1 0 31556 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636968456
transform 1 0 32660 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636968456
transform 1 0 33764 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1
transform 1 0 34868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1
transform 1 0 35420 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636968456
transform 1 0 35604 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636968456
transform 1 0 36708 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636968456
transform 1 0 37812 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1636968456
transform 1 0 38916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1
transform 1 0 40020 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1
transform 1 0 40572 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636968456
transform 1 0 40756 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636968456
transform 1 0 41860 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1636968456
transform 1 0 42964 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1636968456
transform 1 0 44068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1
transform 1 0 45172 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1
transform 1 0 45724 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1636968456
transform 1 0 45908 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1636968456
transform 1 0 47012 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1636968456
transform 1 0 48116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1636968456
transform 1 0 49220 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1
transform 1 0 50324 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1
transform 1 0 50876 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1636968456
transform 1 0 51060 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1636968456
transform 1 0 52164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1636968456
transform 1 0 53268 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1636968456
transform 1 0 54372 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1
transform 1 0 55476 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1
transform 1 0 56028 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1636968456
transform 1 0 56212 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1636968456
transform 1 0 57316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1636968456
transform 1 0 58420 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1636968456
transform 1 0 59524 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1
transform 1 0 60628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1
transform 1 0 61180 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1636968456
transform 1 0 61364 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1636968456
transform 1 0 62468 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1636968456
transform 1 0 63572 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1636968456
transform 1 0 64676 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1
transform 1 0 65780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1
transform 1 0 66332 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1636968456
transform 1 0 66516 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1636968456
transform 1 0 67620 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1636968456
transform 1 0 68724 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1636968456
transform 1 0 69828 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1
transform 1 0 70932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1
transform 1 0 71484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1636968456
transform 1 0 71668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1636968456
transform 1 0 72772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1636968456
transform 1 0 73876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1636968456
transform 1 0 74980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1
transform 1 0 76084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1
transform 1 0 76636 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_813
timestamp 1
transform 1 0 76820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_821
timestamp 1
transform 1 0 77556 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636968456
transform 1 0 2300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636968456
transform 1 0 3404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636968456
transform 1 0 4508 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636968456
transform 1 0 5612 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1
transform 1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636968456
transform 1 0 7268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636968456
transform 1 0 8372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636968456
transform 1 0 9476 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636968456
transform 1 0 10580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1
transform 1 0 11684 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636968456
transform 1 0 12420 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636968456
transform 1 0 13524 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636968456
transform 1 0 14628 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636968456
transform 1 0 15732 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1
transform 1 0 16836 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 17388 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636968456
transform 1 0 17572 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636968456
transform 1 0 18676 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636968456
transform 1 0 19780 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636968456
transform 1 0 20884 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1
transform 1 0 21988 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1
transform 1 0 22540 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636968456
transform 1 0 22724 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636968456
transform 1 0 23828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636968456
transform 1 0 24932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636968456
transform 1 0 26036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1
transform 1 0 27140 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1
transform 1 0 27692 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636968456
transform 1 0 27876 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636968456
transform 1 0 28980 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636968456
transform 1 0 30084 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636968456
transform 1 0 31188 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1
transform 1 0 32292 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1
transform 1 0 32844 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636968456
transform 1 0 33028 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636968456
transform 1 0 34132 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636968456
transform 1 0 35236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636968456
transform 1 0 36340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1
transform 1 0 37444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1
transform 1 0 37996 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636968456
transform 1 0 38180 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636968456
transform 1 0 39284 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636968456
transform 1 0 40388 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636968456
transform 1 0 41492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1
transform 1 0 42596 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1
transform 1 0 43148 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1636968456
transform 1 0 43332 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1636968456
transform 1 0 44436 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1636968456
transform 1 0 45540 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1636968456
transform 1 0 46644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1
transform 1 0 47748 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1
transform 1 0 48300 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1636968456
transform 1 0 48484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1636968456
transform 1 0 49588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1636968456
transform 1 0 50692 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1636968456
transform 1 0 51796 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1
transform 1 0 52900 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1
transform 1 0 53452 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1636968456
transform 1 0 53636 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1636968456
transform 1 0 54740 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1636968456
transform 1 0 55844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1636968456
transform 1 0 56948 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1
transform 1 0 58052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1
transform 1 0 58604 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1636968456
transform 1 0 58788 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1636968456
transform 1 0 59892 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1636968456
transform 1 0 60996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1636968456
transform 1 0 62100 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1
transform 1 0 63204 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1
transform 1 0 63756 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1636968456
transform 1 0 63940 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1636968456
transform 1 0 65044 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1636968456
transform 1 0 66148 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1636968456
transform 1 0 67252 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1
transform 1 0 68356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1
transform 1 0 68908 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1636968456
transform 1 0 69092 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1636968456
transform 1 0 70196 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1636968456
transform 1 0 71300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1636968456
transform 1 0 72404 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1
transform 1 0 73508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1
transform 1 0 74060 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1636968456
transform 1 0 74244 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1636968456
transform 1 0 75348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1636968456
transform 1 0 76452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_821
timestamp 1
transform 1 0 77556 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 3404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 4692 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636968456
transform 1 0 5796 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636968456
transform 1 0 6900 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636968456
transform 1 0 8004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1
transform 1 0 9108 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 9660 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636968456
transform 1 0 9844 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636968456
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636968456
transform 1 0 12052 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636968456
transform 1 0 13156 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1
transform 1 0 14260 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 14812 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636968456
transform 1 0 14996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636968456
transform 1 0 16100 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636968456
transform 1 0 17204 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636968456
transform 1 0 18308 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1
transform 1 0 19412 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1
transform 1 0 19964 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636968456
transform 1 0 20148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636968456
transform 1 0 21252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636968456
transform 1 0 22356 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636968456
transform 1 0 23460 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1
transform 1 0 24564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1
transform 1 0 25116 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636968456
transform 1 0 25300 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636968456
transform 1 0 26404 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636968456
transform 1 0 27508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636968456
transform 1 0 28612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1
transform 1 0 29716 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1
transform 1 0 30268 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636968456
transform 1 0 30452 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636968456
transform 1 0 31556 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636968456
transform 1 0 32660 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636968456
transform 1 0 33764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1
transform 1 0 34868 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1
transform 1 0 35420 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636968456
transform 1 0 35604 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636968456
transform 1 0 36708 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636968456
transform 1 0 37812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1636968456
transform 1 0 38916 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1
transform 1 0 40020 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1
transform 1 0 40572 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636968456
transform 1 0 40756 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636968456
transform 1 0 41860 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636968456
transform 1 0 42964 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1636968456
transform 1 0 44068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1
transform 1 0 45172 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1
transform 1 0 45724 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1636968456
transform 1 0 45908 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1636968456
transform 1 0 47012 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1636968456
transform 1 0 48116 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1636968456
transform 1 0 49220 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1
transform 1 0 50324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1
transform 1 0 50876 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1636968456
transform 1 0 51060 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1636968456
transform 1 0 52164 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1636968456
transform 1 0 53268 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1636968456
transform 1 0 54372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1
transform 1 0 55476 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1
transform 1 0 56028 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1636968456
transform 1 0 56212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1636968456
transform 1 0 57316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1636968456
transform 1 0 58420 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1636968456
transform 1 0 59524 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1
transform 1 0 60628 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1
transform 1 0 61180 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1636968456
transform 1 0 61364 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1636968456
transform 1 0 62468 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1636968456
transform 1 0 63572 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1636968456
transform 1 0 64676 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1
transform 1 0 65780 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1
transform 1 0 66332 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1636968456
transform 1 0 66516 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1636968456
transform 1 0 67620 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1636968456
transform 1 0 68724 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1636968456
transform 1 0 69828 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1
transform 1 0 70932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1
transform 1 0 71484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1636968456
transform 1 0 71668 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1636968456
transform 1 0 72772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1636968456
transform 1 0 73876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1636968456
transform 1 0 74980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1
transform 1 0 76084 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1
transform 1 0 76636 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_813
timestamp 1
transform 1 0 76820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_821
timestamp 1
transform 1 0 77556 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636968456
transform 1 0 2300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636968456
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636968456
transform 1 0 4508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636968456
transform 1 0 5612 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1
transform 1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636968456
transform 1 0 7268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636968456
transform 1 0 8372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636968456
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636968456
transform 1 0 10580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1
transform 1 0 11684 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636968456
transform 1 0 12420 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636968456
transform 1 0 13524 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1636968456
transform 1 0 14628 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1636968456
transform 1 0 15732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1
transform 1 0 16836 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1
transform 1 0 17388 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636968456
transform 1 0 17572 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636968456
transform 1 0 18676 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1636968456
transform 1 0 19780 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1636968456
transform 1 0 20884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1
transform 1 0 21988 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1
transform 1 0 22540 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636968456
transform 1 0 22724 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636968456
transform 1 0 23828 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1636968456
transform 1 0 24932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1636968456
transform 1 0 26036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1
transform 1 0 27140 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1
transform 1 0 27692 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636968456
transform 1 0 27876 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636968456
transform 1 0 28980 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636968456
transform 1 0 30084 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1636968456
transform 1 0 31188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1
transform 1 0 32292 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1
transform 1 0 32844 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636968456
transform 1 0 33028 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1636968456
transform 1 0 34132 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1636968456
transform 1 0 35236 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1636968456
transform 1 0 36340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1
transform 1 0 37444 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1
transform 1 0 37996 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636968456
transform 1 0 38180 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1636968456
transform 1 0 39284 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1636968456
transform 1 0 40388 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1636968456
transform 1 0 41492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1
transform 1 0 42596 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1
transform 1 0 43148 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1636968456
transform 1 0 43332 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1636968456
transform 1 0 44436 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1636968456
transform 1 0 45540 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1636968456
transform 1 0 46644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1
transform 1 0 47748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1
transform 1 0 48300 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1636968456
transform 1 0 48484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1636968456
transform 1 0 49588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1636968456
transform 1 0 50692 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1636968456
transform 1 0 51796 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1
transform 1 0 52900 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1
transform 1 0 53452 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1636968456
transform 1 0 53636 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1636968456
transform 1 0 54740 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1636968456
transform 1 0 55844 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1636968456
transform 1 0 56948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1
transform 1 0 58052 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1
transform 1 0 58604 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1636968456
transform 1 0 58788 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1636968456
transform 1 0 59892 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1636968456
transform 1 0 60996 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1636968456
transform 1 0 62100 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1
transform 1 0 63204 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1
transform 1 0 63756 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1636968456
transform 1 0 63940 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1636968456
transform 1 0 65044 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1636968456
transform 1 0 66148 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1636968456
transform 1 0 67252 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1
transform 1 0 68356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1
transform 1 0 68908 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1636968456
transform 1 0 69092 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1636968456
transform 1 0 70196 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1636968456
transform 1 0 71300 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1636968456
transform 1 0 72404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1
transform 1 0 73508 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1
transform 1 0 74060 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1636968456
transform 1 0 74244 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1636968456
transform 1 0 75348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1636968456
transform 1 0 76452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_821
timestamp 1
transform 1 0 77556 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636968456
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636968456
transform 1 0 3404 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 4508 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636968456
transform 1 0 4692 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636968456
transform 1 0 5796 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636968456
transform 1 0 6900 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636968456
transform 1 0 8004 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1
transform 1 0 9108 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636968456
transform 1 0 9844 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636968456
transform 1 0 10948 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636968456
transform 1 0 12052 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636968456
transform 1 0 13156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1
transform 1 0 14260 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1
transform 1 0 14812 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636968456
transform 1 0 14996 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636968456
transform 1 0 16100 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636968456
transform 1 0 17204 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636968456
transform 1 0 18308 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1
transform 1 0 19412 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636968456
transform 1 0 20148 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1636968456
transform 1 0 21252 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1636968456
transform 1 0 22356 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1636968456
transform 1 0 23460 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1
transform 1 0 24564 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1
transform 1 0 25116 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636968456
transform 1 0 25300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636968456
transform 1 0 26404 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1636968456
transform 1 0 27508 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1636968456
transform 1 0 28612 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1
transform 1 0 29716 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1
transform 1 0 30268 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1636968456
transform 1 0 30452 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1636968456
transform 1 0 31556 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1636968456
transform 1 0 32660 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1636968456
transform 1 0 33764 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1
transform 1 0 34868 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1
transform 1 0 35420 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1636968456
transform 1 0 35604 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1636968456
transform 1 0 36708 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1636968456
transform 1 0 37812 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1636968456
transform 1 0 38916 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1
transform 1 0 40020 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1
transform 1 0 40572 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1636968456
transform 1 0 40756 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1636968456
transform 1 0 41860 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1636968456
transform 1 0 42964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1636968456
transform 1 0 44068 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1
transform 1 0 45172 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1
transform 1 0 45724 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1636968456
transform 1 0 45908 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1636968456
transform 1 0 47012 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1636968456
transform 1 0 48116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1636968456
transform 1 0 49220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1
transform 1 0 50324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1
transform 1 0 50876 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1636968456
transform 1 0 51060 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1636968456
transform 1 0 52164 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1636968456
transform 1 0 53268 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1636968456
transform 1 0 54372 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1
transform 1 0 55476 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1
transform 1 0 56028 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1636968456
transform 1 0 56212 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1636968456
transform 1 0 57316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1636968456
transform 1 0 58420 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1636968456
transform 1 0 59524 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1
transform 1 0 60628 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1
transform 1 0 61180 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1636968456
transform 1 0 61364 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1636968456
transform 1 0 62468 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1636968456
transform 1 0 63572 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1636968456
transform 1 0 64676 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1
transform 1 0 65780 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1
transform 1 0 66332 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1636968456
transform 1 0 66516 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1636968456
transform 1 0 67620 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1636968456
transform 1 0 68724 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1636968456
transform 1 0 69828 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1
transform 1 0 70932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1
transform 1 0 71484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1636968456
transform 1 0 71668 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1636968456
transform 1 0 72772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1636968456
transform 1 0 73876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1636968456
transform 1 0 74980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1
transform 1 0 76084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1
transform 1 0 76636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_813
timestamp 1
transform 1 0 76820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_821
timestamp 1
transform 1 0 77556 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636968456
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636968456
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636968456
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636968456
transform 1 0 5612 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1
transform 1 0 7084 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636968456
transform 1 0 7268 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1636968456
transform 1 0 8372 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1636968456
transform 1 0 9476 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1636968456
transform 1 0 10580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1
transform 1 0 11684 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1
transform 1 0 12236 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636968456
transform 1 0 12420 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1636968456
transform 1 0 13524 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1636968456
transform 1 0 14628 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1636968456
transform 1 0 15732 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1
transform 1 0 16836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1636968456
transform 1 0 17572 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1636968456
transform 1 0 18676 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1636968456
transform 1 0 19780 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1636968456
transform 1 0 20884 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1
transform 1 0 21988 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1
transform 1 0 22540 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636968456
transform 1 0 22724 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636968456
transform 1 0 23828 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1636968456
transform 1 0 24932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1636968456
transform 1 0 26036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1
transform 1 0 27140 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1
transform 1 0 27692 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636968456
transform 1 0 27876 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1636968456
transform 1 0 28980 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1636968456
transform 1 0 30084 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1636968456
transform 1 0 31188 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1
transform 1 0 32292 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1
transform 1 0 32844 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1636968456
transform 1 0 33028 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1636968456
transform 1 0 34132 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1636968456
transform 1 0 35236 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1636968456
transform 1 0 36340 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1
transform 1 0 37444 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1
transform 1 0 37996 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1636968456
transform 1 0 38180 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1636968456
transform 1 0 39284 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1636968456
transform 1 0 40388 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1636968456
transform 1 0 41492 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1
transform 1 0 42596 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1
transform 1 0 43148 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1636968456
transform 1 0 43332 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1636968456
transform 1 0 44436 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1636968456
transform 1 0 45540 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1636968456
transform 1 0 46644 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1
transform 1 0 47748 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1
transform 1 0 48300 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1636968456
transform 1 0 48484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1636968456
transform 1 0 49588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1636968456
transform 1 0 50692 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1636968456
transform 1 0 51796 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1
transform 1 0 52900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1
transform 1 0 53452 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1636968456
transform 1 0 53636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1636968456
transform 1 0 54740 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1636968456
transform 1 0 55844 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1636968456
transform 1 0 56948 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1
transform 1 0 58052 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1
transform 1 0 58604 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1636968456
transform 1 0 58788 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1636968456
transform 1 0 59892 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1636968456
transform 1 0 60996 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1636968456
transform 1 0 62100 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1
transform 1 0 63204 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1
transform 1 0 63756 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1636968456
transform 1 0 63940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1636968456
transform 1 0 65044 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1636968456
transform 1 0 66148 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1636968456
transform 1 0 67252 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1
transform 1 0 68356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1
transform 1 0 68908 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1636968456
transform 1 0 69092 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1636968456
transform 1 0 70196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1636968456
transform 1 0 71300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1636968456
transform 1 0 72404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1
transform 1 0 73508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1
transform 1 0 74060 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1636968456
transform 1 0 74244 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1636968456
transform 1 0 75348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1636968456
transform 1 0 76452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_821
timestamp 1
transform 1 0 77556 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636968456
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636968456
transform 1 0 3404 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636968456
transform 1 0 4692 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636968456
transform 1 0 5796 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636968456
transform 1 0 6900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1636968456
transform 1 0 8004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1
transform 1 0 9108 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1636968456
transform 1 0 9844 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1636968456
transform 1 0 10948 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1636968456
transform 1 0 12052 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1636968456
transform 1 0 13156 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1
transform 1 0 14260 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636968456
transform 1 0 14996 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636968456
transform 1 0 16100 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1636968456
transform 1 0 17204 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1636968456
transform 1 0 18308 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1
transform 1 0 19412 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1
transform 1 0 19964 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1636968456
transform 1 0 20148 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1636968456
transform 1 0 21252 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1636968456
transform 1 0 22356 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1636968456
transform 1 0 23460 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1
transform 1 0 24564 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1
transform 1 0 25116 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1636968456
transform 1 0 25300 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1636968456
transform 1 0 26404 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1636968456
transform 1 0 27508 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1636968456
transform 1 0 28612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1
transform 1 0 29716 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1
transform 1 0 30268 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1636968456
transform 1 0 30452 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1636968456
transform 1 0 31556 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1636968456
transform 1 0 32660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1636968456
transform 1 0 33764 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1
transform 1 0 34868 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1
transform 1 0 35420 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1636968456
transform 1 0 35604 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1636968456
transform 1 0 36708 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1636968456
transform 1 0 37812 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1636968456
transform 1 0 38916 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1
transform 1 0 40020 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1
transform 1 0 40572 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1636968456
transform 1 0 40756 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1636968456
transform 1 0 41860 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1636968456
transform 1 0 42964 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1636968456
transform 1 0 44068 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1
transform 1 0 45172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1
transform 1 0 45724 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1636968456
transform 1 0 45908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1636968456
transform 1 0 47012 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1636968456
transform 1 0 48116 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1636968456
transform 1 0 49220 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1
transform 1 0 50324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1
transform 1 0 50876 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1636968456
transform 1 0 51060 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1636968456
transform 1 0 52164 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1636968456
transform 1 0 53268 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1636968456
transform 1 0 54372 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1
transform 1 0 55476 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1
transform 1 0 56028 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1636968456
transform 1 0 56212 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1636968456
transform 1 0 57316 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1636968456
transform 1 0 58420 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1636968456
transform 1 0 59524 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1
transform 1 0 60628 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1
transform 1 0 61180 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1636968456
transform 1 0 61364 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1636968456
transform 1 0 62468 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1636968456
transform 1 0 63572 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1636968456
transform 1 0 64676 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1
transform 1 0 65780 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1
transform 1 0 66332 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1636968456
transform 1 0 66516 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1636968456
transform 1 0 67620 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_725
timestamp 1636968456
transform 1 0 68724 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_737
timestamp 1636968456
transform 1 0 69828 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1
transform 1 0 70932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1
transform 1 0 71484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1636968456
transform 1 0 71668 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1636968456
transform 1 0 72772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1636968456
transform 1 0 73876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1636968456
transform 1 0 74980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1
transform 1 0 76084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1
transform 1 0 76636 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_813
timestamp 1
transform 1 0 76820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_821
timestamp 1
transform 1 0 77556 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 2300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636968456
transform 1 0 3404 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636968456
transform 1 0 4508 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636968456
transform 1 0 5612 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636968456
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636968456
transform 1 0 8372 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1636968456
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1636968456
transform 1 0 10580 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1
transform 1 0 11684 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1636968456
transform 1 0 12420 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1636968456
transform 1 0 13524 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1636968456
transform 1 0 14628 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1636968456
transform 1 0 15732 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1
transform 1 0 16836 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636968456
transform 1 0 17572 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1636968456
transform 1 0 18676 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1636968456
transform 1 0 19780 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1636968456
transform 1 0 20884 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1
transform 1 0 21988 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1
transform 1 0 22540 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1636968456
transform 1 0 22724 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1636968456
transform 1 0 23828 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1636968456
transform 1 0 24932 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1636968456
transform 1 0 26036 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1
transform 1 0 27140 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1
transform 1 0 27692 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1636968456
transform 1 0 27876 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1636968456
transform 1 0 28980 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1636968456
transform 1 0 30084 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1636968456
transform 1 0 31188 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1
transform 1 0 32292 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1
transform 1 0 32844 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1636968456
transform 1 0 33028 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1636968456
transform 1 0 34132 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1636968456
transform 1 0 35236 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1636968456
transform 1 0 36340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1
transform 1 0 37444 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1
transform 1 0 37996 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1636968456
transform 1 0 38180 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1636968456
transform 1 0 39284 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1636968456
transform 1 0 40388 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1636968456
transform 1 0 41492 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1
transform 1 0 42596 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1
transform 1 0 43148 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1636968456
transform 1 0 43332 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1636968456
transform 1 0 44436 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1636968456
transform 1 0 45540 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1636968456
transform 1 0 46644 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1
transform 1 0 47748 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1
transform 1 0 48300 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1636968456
transform 1 0 48484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1636968456
transform 1 0 49588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1636968456
transform 1 0 50692 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1636968456
transform 1 0 51796 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1
transform 1 0 52900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1
transform 1 0 53452 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1636968456
transform 1 0 53636 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1636968456
transform 1 0 54740 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1636968456
transform 1 0 55844 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1636968456
transform 1 0 56948 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1
transform 1 0 58052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1
transform 1 0 58604 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1636968456
transform 1 0 58788 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1636968456
transform 1 0 59892 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1636968456
transform 1 0 60996 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1636968456
transform 1 0 62100 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1
transform 1 0 63204 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1
transform 1 0 63756 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1636968456
transform 1 0 63940 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1636968456
transform 1 0 65044 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1636968456
transform 1 0 66148 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1636968456
transform 1 0 67252 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1
transform 1 0 68356 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1
transform 1 0 68908 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1636968456
transform 1 0 69092 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1636968456
transform 1 0 70196 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_753
timestamp 1636968456
transform 1 0 71300 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_765
timestamp 1636968456
transform 1 0 72404 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1
transform 1 0 73508 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1
transform 1 0 74060 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1636968456
transform 1 0 74244 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1636968456
transform 1 0 75348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_809
timestamp 1636968456
transform 1 0 76452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_821
timestamp 1
transform 1 0 77556 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636968456
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636968456
transform 1 0 3404 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636968456
transform 1 0 4692 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636968456
transform 1 0 5796 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636968456
transform 1 0 6900 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1636968456
transform 1 0 8004 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1
transform 1 0 9108 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636968456
transform 1 0 9844 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636968456
transform 1 0 10948 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1636968456
transform 1 0 12052 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1636968456
transform 1 0 13156 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1
transform 1 0 14260 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636968456
transform 1 0 14996 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1636968456
transform 1 0 16100 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1636968456
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1636968456
transform 1 0 18308 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1
transform 1 0 19412 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1636968456
transform 1 0 20148 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1636968456
transform 1 0 21252 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1636968456
transform 1 0 22356 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1636968456
transform 1 0 23460 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1
transform 1 0 24564 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1
transform 1 0 25116 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1636968456
transform 1 0 25300 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1636968456
transform 1 0 26404 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1636968456
transform 1 0 27508 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1636968456
transform 1 0 28612 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1
transform 1 0 29716 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1
transform 1 0 30268 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1636968456
transform 1 0 30452 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1636968456
transform 1 0 31556 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1636968456
transform 1 0 32660 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1636968456
transform 1 0 33764 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1
transform 1 0 34868 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1
transform 1 0 35420 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1636968456
transform 1 0 35604 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1636968456
transform 1 0 36708 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1636968456
transform 1 0 37812 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1636968456
transform 1 0 38916 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1
transform 1 0 40020 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1
transform 1 0 40572 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1636968456
transform 1 0 40756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1636968456
transform 1 0 41860 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1636968456
transform 1 0 42964 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1636968456
transform 1 0 44068 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1
transform 1 0 45172 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1
transform 1 0 45724 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1636968456
transform 1 0 45908 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1636968456
transform 1 0 47012 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1636968456
transform 1 0 48116 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1636968456
transform 1 0 49220 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1
transform 1 0 50324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1
transform 1 0 50876 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1636968456
transform 1 0 51060 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1636968456
transform 1 0 52164 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1636968456
transform 1 0 53268 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1636968456
transform 1 0 54372 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1
transform 1 0 55476 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1
transform 1 0 56028 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1636968456
transform 1 0 56212 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1636968456
transform 1 0 57316 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1636968456
transform 1 0 58420 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1636968456
transform 1 0 59524 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1
transform 1 0 60628 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1
transform 1 0 61180 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1636968456
transform 1 0 61364 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1636968456
transform 1 0 62468 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1636968456
transform 1 0 63572 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1636968456
transform 1 0 64676 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1
transform 1 0 65780 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1
transform 1 0 66332 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1636968456
transform 1 0 66516 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1636968456
transform 1 0 67620 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_725
timestamp 1636968456
transform 1 0 68724 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_737
timestamp 1636968456
transform 1 0 69828 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1
transform 1 0 70932 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1
transform 1 0 71484 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_757
timestamp 1636968456
transform 1 0 71668 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_769
timestamp 1636968456
transform 1 0 72772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_781
timestamp 1636968456
transform 1 0 73876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_793
timestamp 1636968456
transform 1 0 74980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1
transform 1 0 76084 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1
transform 1 0 76636 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_813
timestamp 1
transform 1 0 76820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_821
timestamp 1
transform 1 0 77556 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636968456
transform 1 0 2300 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636968456
transform 1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636968456
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636968456
transform 1 0 5612 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636968456
transform 1 0 7268 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1636968456
transform 1 0 8372 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1636968456
transform 1 0 9476 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1636968456
transform 1 0 10580 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1
transform 1 0 11684 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1
transform 1 0 12236 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1636968456
transform 1 0 12420 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1636968456
transform 1 0 13524 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1636968456
transform 1 0 14628 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1636968456
transform 1 0 15732 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1
transform 1 0 16836 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636968456
transform 1 0 17572 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1636968456
transform 1 0 18676 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1636968456
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1636968456
transform 1 0 20884 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1
transform 1 0 21988 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1
transform 1 0 22540 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1636968456
transform 1 0 22724 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1636968456
transform 1 0 23828 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1636968456
transform 1 0 24932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1636968456
transform 1 0 26036 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1
transform 1 0 27140 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1
transform 1 0 27692 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1636968456
transform 1 0 27876 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1636968456
transform 1 0 28980 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1636968456
transform 1 0 30084 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1636968456
transform 1 0 31188 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1
transform 1 0 32292 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1
transform 1 0 32844 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1636968456
transform 1 0 33028 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1636968456
transform 1 0 34132 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1636968456
transform 1 0 35236 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1636968456
transform 1 0 36340 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1
transform 1 0 37444 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1
transform 1 0 37996 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1636968456
transform 1 0 38180 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1636968456
transform 1 0 39284 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1636968456
transform 1 0 40388 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1636968456
transform 1 0 41492 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1
transform 1 0 42596 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1
transform 1 0 43148 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1636968456
transform 1 0 43332 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1636968456
transform 1 0 44436 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1636968456
transform 1 0 45540 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1636968456
transform 1 0 46644 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1
transform 1 0 47748 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1
transform 1 0 48300 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1636968456
transform 1 0 48484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1636968456
transform 1 0 49588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1636968456
transform 1 0 50692 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1636968456
transform 1 0 51796 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1
transform 1 0 52900 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1
transform 1 0 53452 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1636968456
transform 1 0 53636 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1636968456
transform 1 0 54740 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1636968456
transform 1 0 55844 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1636968456
transform 1 0 56948 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1
transform 1 0 58052 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1
transform 1 0 58604 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1636968456
transform 1 0 58788 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1636968456
transform 1 0 59892 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1636968456
transform 1 0 60996 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1636968456
transform 1 0 62100 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1
transform 1 0 63204 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1
transform 1 0 63756 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1636968456
transform 1 0 63940 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1636968456
transform 1 0 65044 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1636968456
transform 1 0 66148 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1636968456
transform 1 0 67252 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1
transform 1 0 68356 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1
transform 1 0 68908 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_729
timestamp 1636968456
transform 1 0 69092 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_741
timestamp 1636968456
transform 1 0 70196 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_753
timestamp 1636968456
transform 1 0 71300 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_765
timestamp 1636968456
transform 1 0 72404 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1
transform 1 0 73508 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1
transform 1 0 74060 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_785
timestamp 1636968456
transform 1 0 74244 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_797
timestamp 1636968456
transform 1 0 75348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_809
timestamp 1636968456
transform 1 0 76452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_821
timestamp 1
transform 1 0 77556 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636968456
transform 1 0 2300 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636968456
transform 1 0 3404 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636968456
transform 1 0 4692 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636968456
transform 1 0 5796 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636968456
transform 1 0 6900 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1636968456
transform 1 0 8004 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1
transform 1 0 9108 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1
transform 1 0 9660 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636968456
transform 1 0 9844 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1636968456
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1636968456
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1636968456
transform 1 0 13156 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1
transform 1 0 14260 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1
transform 1 0 14812 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636968456
transform 1 0 14996 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1636968456
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1636968456
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1636968456
transform 1 0 18308 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1
transform 1 0 19412 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1
transform 1 0 19964 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1636968456
transform 1 0 20148 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1636968456
transform 1 0 21252 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1636968456
transform 1 0 22356 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1636968456
transform 1 0 23460 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1
transform 1 0 24564 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1
transform 1 0 25116 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1636968456
transform 1 0 25300 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1636968456
transform 1 0 26404 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1636968456
transform 1 0 27508 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1636968456
transform 1 0 28612 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1
transform 1 0 29716 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1
transform 1 0 30268 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1636968456
transform 1 0 30452 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1636968456
transform 1 0 31556 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1636968456
transform 1 0 32660 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1636968456
transform 1 0 33764 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1
transform 1 0 34868 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1
transform 1 0 35420 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1636968456
transform 1 0 35604 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1636968456
transform 1 0 36708 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1636968456
transform 1 0 37812 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1636968456
transform 1 0 38916 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1
transform 1 0 40020 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1
transform 1 0 40572 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1636968456
transform 1 0 40756 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1636968456
transform 1 0 41860 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1636968456
transform 1 0 42964 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1636968456
transform 1 0 44068 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1
transform 1 0 45172 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1
transform 1 0 45724 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1636968456
transform 1 0 45908 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1636968456
transform 1 0 47012 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1636968456
transform 1 0 48116 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1636968456
transform 1 0 49220 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1
transform 1 0 50324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1
transform 1 0 50876 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1636968456
transform 1 0 51060 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1636968456
transform 1 0 52164 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1636968456
transform 1 0 53268 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1636968456
transform 1 0 54372 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1
transform 1 0 55476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1
transform 1 0 56028 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1636968456
transform 1 0 56212 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1636968456
transform 1 0 57316 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1636968456
transform 1 0 58420 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1636968456
transform 1 0 59524 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1
transform 1 0 60628 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1
transform 1 0 61180 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1636968456
transform 1 0 61364 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1636968456
transform 1 0 62468 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1636968456
transform 1 0 63572 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1636968456
transform 1 0 64676 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1
transform 1 0 65780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1
transform 1 0 66332 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1636968456
transform 1 0 66516 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1636968456
transform 1 0 67620 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_725
timestamp 1636968456
transform 1 0 68724 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_737
timestamp 1636968456
transform 1 0 69828 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1
transform 1 0 70932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1
transform 1 0 71484 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_757
timestamp 1636968456
transform 1 0 71668 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_769
timestamp 1636968456
transform 1 0 72772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_781
timestamp 1636968456
transform 1 0 73876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_793
timestamp 1636968456
transform 1 0 74980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1
transform 1 0 76084 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1
transform 1 0 76636 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_813
timestamp 1
transform 1 0 76820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_821
timestamp 1
transform 1 0 77556 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636968456
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636968456
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636968456
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1636968456
transform 1 0 5612 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1
transform 1 0 6716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636968456
transform 1 0 7268 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636968456
transform 1 0 8372 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1636968456
transform 1 0 9476 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1636968456
transform 1 0 10580 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1
transform 1 0 11684 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636968456
transform 1 0 12420 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1636968456
transform 1 0 13524 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1636968456
transform 1 0 14628 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1636968456
transform 1 0 15732 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1
transform 1 0 16836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1
transform 1 0 17388 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636968456
transform 1 0 17572 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1636968456
transform 1 0 18676 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1636968456
transform 1 0 19780 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1636968456
transform 1 0 20884 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1
transform 1 0 21988 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1
transform 1 0 22540 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1636968456
transform 1 0 22724 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1636968456
transform 1 0 23828 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1636968456
transform 1 0 24932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1636968456
transform 1 0 26036 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1
transform 1 0 27140 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1
transform 1 0 27692 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1636968456
transform 1 0 27876 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1636968456
transform 1 0 28980 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1636968456
transform 1 0 30084 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1636968456
transform 1 0 31188 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1
transform 1 0 32292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1
transform 1 0 32844 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1636968456
transform 1 0 33028 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1636968456
transform 1 0 34132 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1636968456
transform 1 0 35236 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1636968456
transform 1 0 36340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1
transform 1 0 37444 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1
transform 1 0 37996 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1636968456
transform 1 0 38180 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1636968456
transform 1 0 39284 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1636968456
transform 1 0 40388 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1636968456
transform 1 0 41492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1
transform 1 0 42596 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1
transform 1 0 43148 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1636968456
transform 1 0 43332 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1636968456
transform 1 0 44436 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1636968456
transform 1 0 45540 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1636968456
transform 1 0 46644 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1
transform 1 0 47748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1
transform 1 0 48300 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1636968456
transform 1 0 48484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1636968456
transform 1 0 49588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1636968456
transform 1 0 50692 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1636968456
transform 1 0 51796 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1
transform 1 0 52900 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1
transform 1 0 53452 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1636968456
transform 1 0 53636 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1636968456
transform 1 0 54740 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1636968456
transform 1 0 55844 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1636968456
transform 1 0 56948 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1
transform 1 0 58052 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1
transform 1 0 58604 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1636968456
transform 1 0 58788 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1636968456
transform 1 0 59892 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1636968456
transform 1 0 60996 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1636968456
transform 1 0 62100 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1
transform 1 0 63204 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1
transform 1 0 63756 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1636968456
transform 1 0 63940 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1636968456
transform 1 0 65044 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1636968456
transform 1 0 66148 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1636968456
transform 1 0 67252 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1
transform 1 0 68356 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1
transform 1 0 68908 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_729
timestamp 1636968456
transform 1 0 69092 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_741
timestamp 1636968456
transform 1 0 70196 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_753
timestamp 1636968456
transform 1 0 71300 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_765
timestamp 1636968456
transform 1 0 72404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1
transform 1 0 73508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1
transform 1 0 74060 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_785
timestamp 1636968456
transform 1 0 74244 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_797
timestamp 1636968456
transform 1 0 75348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_809
timestamp 1636968456
transform 1 0 76452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_821
timestamp 1
transform 1 0 77556 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636968456
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636968456
transform 1 0 3404 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636968456
transform 1 0 4692 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636968456
transform 1 0 5796 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636968456
transform 1 0 6900 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1636968456
transform 1 0 8004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1
transform 1 0 9108 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636968456
transform 1 0 9844 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636968456
transform 1 0 10948 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1636968456
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1636968456
transform 1 0 13156 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1
transform 1 0 14260 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636968456
transform 1 0 14996 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636968456
transform 1 0 16100 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636968456
transform 1 0 17204 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1636968456
transform 1 0 18308 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1
transform 1 0 19412 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1636968456
transform 1 0 20148 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1636968456
transform 1 0 21252 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1636968456
transform 1 0 22356 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1636968456
transform 1 0 23460 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1
transform 1 0 24564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1
transform 1 0 25116 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1636968456
transform 1 0 25300 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1636968456
transform 1 0 26404 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1636968456
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1636968456
transform 1 0 28612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1
transform 1 0 29716 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1
transform 1 0 30268 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1636968456
transform 1 0 30452 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1636968456
transform 1 0 31556 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1636968456
transform 1 0 32660 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1636968456
transform 1 0 33764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1
transform 1 0 34868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1
transform 1 0 35420 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1636968456
transform 1 0 35604 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1636968456
transform 1 0 36708 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1636968456
transform 1 0 37812 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1636968456
transform 1 0 38916 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1
transform 1 0 40020 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1
transform 1 0 40572 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1636968456
transform 1 0 40756 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1636968456
transform 1 0 41860 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1636968456
transform 1 0 42964 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1636968456
transform 1 0 44068 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1
transform 1 0 45172 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1
transform 1 0 45724 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1636968456
transform 1 0 45908 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1636968456
transform 1 0 47012 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1636968456
transform 1 0 48116 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1636968456
transform 1 0 49220 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1
transform 1 0 50324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1
transform 1 0 50876 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1636968456
transform 1 0 51060 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1636968456
transform 1 0 52164 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1636968456
transform 1 0 53268 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1636968456
transform 1 0 54372 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1
transform 1 0 55476 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1
transform 1 0 56028 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1636968456
transform 1 0 56212 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1636968456
transform 1 0 57316 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1636968456
transform 1 0 58420 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1636968456
transform 1 0 59524 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1
transform 1 0 60628 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1
transform 1 0 61180 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1636968456
transform 1 0 61364 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1636968456
transform 1 0 62468 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1636968456
transform 1 0 63572 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1636968456
transform 1 0 64676 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1
transform 1 0 65780 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1
transform 1 0 66332 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1636968456
transform 1 0 66516 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1636968456
transform 1 0 67620 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_725
timestamp 1636968456
transform 1 0 68724 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_737
timestamp 1636968456
transform 1 0 69828 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 1
transform 1 0 70932 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1
transform 1 0 71484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_757
timestamp 1636968456
transform 1 0 71668 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_769
timestamp 1636968456
transform 1 0 72772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_781
timestamp 1636968456
transform 1 0 73876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_793
timestamp 1636968456
transform 1 0 74980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_805
timestamp 1
transform 1 0 76084 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 1
transform 1 0 76636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_813
timestamp 1
transform 1 0 76820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_821
timestamp 1
transform 1 0 77556 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636968456
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636968456
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636968456
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636968456
transform 1 0 5612 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1
transform 1 0 6716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636968456
transform 1 0 7268 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636968456
transform 1 0 8372 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1636968456
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1636968456
transform 1 0 10580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1
transform 1 0 11684 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636968456
transform 1 0 12420 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636968456
transform 1 0 13524 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1636968456
transform 1 0 14628 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1636968456
transform 1 0 15732 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1
transform 1 0 16836 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1
transform 1 0 17388 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636968456
transform 1 0 17572 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1636968456
transform 1 0 18676 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1636968456
transform 1 0 19780 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1636968456
transform 1 0 20884 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1
transform 1 0 21988 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1
transform 1 0 22540 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636968456
transform 1 0 22724 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1636968456
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1636968456
transform 1 0 24932 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1636968456
transform 1 0 26036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1
transform 1 0 27140 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1
transform 1 0 27692 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1636968456
transform 1 0 27876 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1636968456
transform 1 0 28980 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1636968456
transform 1 0 30084 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1636968456
transform 1 0 31188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1
transform 1 0 32292 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1
transform 1 0 32844 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1636968456
transform 1 0 33028 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1636968456
transform 1 0 34132 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1636968456
transform 1 0 35236 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1636968456
transform 1 0 36340 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1
transform 1 0 37444 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1636968456
transform 1 0 38180 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1636968456
transform 1 0 39284 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1636968456
transform 1 0 40388 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1636968456
transform 1 0 41492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1
transform 1 0 42596 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1
transform 1 0 43148 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1636968456
transform 1 0 43332 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1636968456
transform 1 0 44436 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1636968456
transform 1 0 45540 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1636968456
transform 1 0 46644 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1
transform 1 0 47748 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1
transform 1 0 48300 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1636968456
transform 1 0 48484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1636968456
transform 1 0 49588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1636968456
transform 1 0 50692 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1636968456
transform 1 0 51796 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1
transform 1 0 52900 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1
transform 1 0 53452 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1636968456
transform 1 0 53636 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1636968456
transform 1 0 54740 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1636968456
transform 1 0 55844 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1636968456
transform 1 0 56948 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1
transform 1 0 58052 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1
transform 1 0 58604 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1636968456
transform 1 0 58788 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1636968456
transform 1 0 59892 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1636968456
transform 1 0 60996 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1636968456
transform 1 0 62100 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1
transform 1 0 63204 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1
transform 1 0 63756 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1636968456
transform 1 0 63940 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1636968456
transform 1 0 65044 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1636968456
transform 1 0 66148 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1636968456
transform 1 0 67252 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1
transform 1 0 68356 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1
transform 1 0 68908 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_729
timestamp 1636968456
transform 1 0 69092 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_741
timestamp 1636968456
transform 1 0 70196 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_753
timestamp 1636968456
transform 1 0 71300 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_765
timestamp 1636968456
transform 1 0 72404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 1
transform 1 0 73508 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1
transform 1 0 74060 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_785
timestamp 1636968456
transform 1 0 74244 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_797
timestamp 1636968456
transform 1 0 75348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_809
timestamp 1636968456
transform 1 0 76452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_821
timestamp 1
transform 1 0 77556 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636968456
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636968456
transform 1 0 3404 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636968456
transform 1 0 4692 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636968456
transform 1 0 5796 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636968456
transform 1 0 6900 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1636968456
transform 1 0 8004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1
transform 1 0 9108 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1
transform 1 0 9660 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636968456
transform 1 0 9844 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636968456
transform 1 0 10948 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636968456
transform 1 0 12052 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1636968456
transform 1 0 13156 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1
transform 1 0 14260 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1
transform 1 0 14812 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636968456
transform 1 0 14996 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1636968456
transform 1 0 16100 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1636968456
transform 1 0 17204 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1636968456
transform 1 0 18308 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1
transform 1 0 19412 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1
transform 1 0 19964 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636968456
transform 1 0 20148 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1636968456
transform 1 0 21252 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1636968456
transform 1 0 22356 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1636968456
transform 1 0 23460 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1
transform 1 0 24564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1
transform 1 0 25116 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1636968456
transform 1 0 25300 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1636968456
transform 1 0 26404 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1636968456
transform 1 0 27508 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1636968456
transform 1 0 28612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1
transform 1 0 29716 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1
transform 1 0 30268 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1636968456
transform 1 0 30452 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1636968456
transform 1 0 31556 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1636968456
transform 1 0 32660 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1636968456
transform 1 0 33764 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1
transform 1 0 34868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1
transform 1 0 35420 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1636968456
transform 1 0 35604 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1636968456
transform 1 0 36708 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1636968456
transform 1 0 37812 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1636968456
transform 1 0 38916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1
transform 1 0 40020 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1
transform 1 0 40572 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1636968456
transform 1 0 40756 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1636968456
transform 1 0 41860 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1636968456
transform 1 0 42964 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1636968456
transform 1 0 44068 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1
transform 1 0 45172 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1
transform 1 0 45724 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1636968456
transform 1 0 45908 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1636968456
transform 1 0 47012 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1636968456
transform 1 0 48116 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1636968456
transform 1 0 49220 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1
transform 1 0 50324 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1
transform 1 0 50876 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1636968456
transform 1 0 51060 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1636968456
transform 1 0 52164 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1636968456
transform 1 0 53268 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1636968456
transform 1 0 54372 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1
transform 1 0 55476 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1
transform 1 0 56028 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1636968456
transform 1 0 56212 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1636968456
transform 1 0 57316 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1636968456
transform 1 0 58420 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1636968456
transform 1 0 59524 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1
transform 1 0 60628 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1
transform 1 0 61180 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1636968456
transform 1 0 61364 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1636968456
transform 1 0 62468 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1636968456
transform 1 0 63572 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1636968456
transform 1 0 64676 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1
transform 1 0 65780 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1
transform 1 0 66332 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1636968456
transform 1 0 66516 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1636968456
transform 1 0 67620 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_725
timestamp 1636968456
transform 1 0 68724 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_737
timestamp 1636968456
transform 1 0 69828 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_749
timestamp 1
transform 1 0 70932 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_755
timestamp 1
transform 1 0 71484 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_757
timestamp 1636968456
transform 1 0 71668 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_769
timestamp 1636968456
transform 1 0 72772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_781
timestamp 1636968456
transform 1 0 73876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_793
timestamp 1636968456
transform 1 0 74980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_805
timestamp 1
transform 1 0 76084 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_811
timestamp 1
transform 1 0 76636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_813
timestamp 1
transform 1 0 76820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_821
timestamp 1
transform 1 0 77556 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636968456
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636968456
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636968456
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636968456
transform 1 0 5612 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1
transform 1 0 6716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636968456
transform 1 0 7268 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1636968456
transform 1 0 8372 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1636968456
transform 1 0 9476 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1636968456
transform 1 0 10580 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1
transform 1 0 11684 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1636968456
transform 1 0 12420 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1636968456
transform 1 0 13524 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1636968456
transform 1 0 14628 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1636968456
transform 1 0 15732 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1
transform 1 0 16836 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1
transform 1 0 17388 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1636968456
transform 1 0 17572 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1636968456
transform 1 0 18676 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1636968456
transform 1 0 19780 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1636968456
transform 1 0 20884 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1
transform 1 0 21988 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1
transform 1 0 22540 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1636968456
transform 1 0 22724 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1636968456
transform 1 0 23828 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1636968456
transform 1 0 24932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1636968456
transform 1 0 26036 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1
transform 1 0 27140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1
transform 1 0 27692 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1636968456
transform 1 0 27876 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1636968456
transform 1 0 28980 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1636968456
transform 1 0 30084 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1636968456
transform 1 0 31188 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1
transform 1 0 32292 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1
transform 1 0 32844 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1636968456
transform 1 0 33028 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1636968456
transform 1 0 34132 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1636968456
transform 1 0 35236 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1636968456
transform 1 0 36340 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1
transform 1 0 37444 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1
transform 1 0 37996 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1636968456
transform 1 0 38180 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1636968456
transform 1 0 39284 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1636968456
transform 1 0 40388 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1636968456
transform 1 0 41492 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1
transform 1 0 42596 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1
transform 1 0 43148 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1636968456
transform 1 0 43332 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1636968456
transform 1 0 44436 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1636968456
transform 1 0 45540 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1636968456
transform 1 0 46644 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1
transform 1 0 47748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1
transform 1 0 48300 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1636968456
transform 1 0 48484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1636968456
transform 1 0 49588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1636968456
transform 1 0 50692 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1636968456
transform 1 0 51796 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1
transform 1 0 52900 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1
transform 1 0 53452 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1636968456
transform 1 0 53636 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1636968456
transform 1 0 54740 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1636968456
transform 1 0 55844 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1636968456
transform 1 0 56948 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1
transform 1 0 58052 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1
transform 1 0 58604 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1636968456
transform 1 0 58788 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1636968456
transform 1 0 59892 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1636968456
transform 1 0 60996 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1636968456
transform 1 0 62100 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1
transform 1 0 63204 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1
transform 1 0 63756 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1636968456
transform 1 0 63940 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1636968456
transform 1 0 65044 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1636968456
transform 1 0 66148 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1636968456
transform 1 0 67252 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1
transform 1 0 68356 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1
transform 1 0 68908 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_729
timestamp 1636968456
transform 1 0 69092 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_741
timestamp 1636968456
transform 1 0 70196 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_753
timestamp 1636968456
transform 1 0 71300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_765
timestamp 1636968456
transform 1 0 72404 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_777
timestamp 1
transform 1 0 73508 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 1
transform 1 0 74060 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_785
timestamp 1636968456
transform 1 0 74244 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_797
timestamp 1636968456
transform 1 0 75348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_809
timestamp 1636968456
transform 1 0 76452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_821
timestamp 1
transform 1 0 77556 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636968456
transform 1 0 2300 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636968456
transform 1 0 3404 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1
transform 1 0 4508 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636968456
transform 1 0 4692 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636968456
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636968456
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1636968456
transform 1 0 8004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1
transform 1 0 9108 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636968456
transform 1 0 9844 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1636968456
transform 1 0 10948 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1636968456
transform 1 0 12052 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1636968456
transform 1 0 13156 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1
transform 1 0 14260 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636968456
transform 1 0 14996 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1636968456
transform 1 0 16100 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1636968456
transform 1 0 17204 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1636968456
transform 1 0 18308 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1
transform 1 0 19412 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1
transform 1 0 19964 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636968456
transform 1 0 20148 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1636968456
transform 1 0 21252 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1636968456
transform 1 0 22356 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1636968456
transform 1 0 23460 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1
transform 1 0 24564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1
transform 1 0 25116 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1636968456
transform 1 0 25300 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1636968456
transform 1 0 26404 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1636968456
transform 1 0 27508 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1636968456
transform 1 0 28612 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1
transform 1 0 29716 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1
transform 1 0 30268 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1636968456
transform 1 0 30452 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1636968456
transform 1 0 31556 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1636968456
transform 1 0 32660 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1636968456
transform 1 0 33764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1
transform 1 0 34868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1
transform 1 0 35420 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1636968456
transform 1 0 35604 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1636968456
transform 1 0 36708 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1636968456
transform 1 0 37812 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1636968456
transform 1 0 38916 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1
transform 1 0 40020 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1
transform 1 0 40572 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1636968456
transform 1 0 40756 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1636968456
transform 1 0 41860 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1636968456
transform 1 0 42964 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1636968456
transform 1 0 44068 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1
transform 1 0 45172 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1
transform 1 0 45724 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1636968456
transform 1 0 45908 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1636968456
transform 1 0 47012 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1636968456
transform 1 0 48116 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1636968456
transform 1 0 49220 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1
transform 1 0 50324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1
transform 1 0 50876 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1636968456
transform 1 0 51060 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1636968456
transform 1 0 52164 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1636968456
transform 1 0 53268 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1636968456
transform 1 0 54372 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1
transform 1 0 55476 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1
transform 1 0 56028 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1636968456
transform 1 0 56212 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1636968456
transform 1 0 57316 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1636968456
transform 1 0 58420 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1636968456
transform 1 0 59524 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1
transform 1 0 60628 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1
transform 1 0 61180 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1636968456
transform 1 0 61364 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1636968456
transform 1 0 62468 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1636968456
transform 1 0 63572 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1636968456
transform 1 0 64676 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1
transform 1 0 65780 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1
transform 1 0 66332 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1636968456
transform 1 0 66516 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1636968456
transform 1 0 67620 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_725
timestamp 1636968456
transform 1 0 68724 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_737
timestamp 1636968456
transform 1 0 69828 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_749
timestamp 1
transform 1 0 70932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_755
timestamp 1
transform 1 0 71484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_757
timestamp 1636968456
transform 1 0 71668 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_769
timestamp 1636968456
transform 1 0 72772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_781
timestamp 1636968456
transform 1 0 73876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_793
timestamp 1636968456
transform 1 0 74980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_805
timestamp 1
transform 1 0 76084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_811
timestamp 1
transform 1 0 76636 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_813
timestamp 1
transform 1 0 76820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_821
timestamp 1
transform 1 0 77556 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636968456
transform 1 0 2300 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636968456
transform 1 0 3404 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636968456
transform 1 0 4508 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636968456
transform 1 0 5612 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1
transform 1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636968456
transform 1 0 7268 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1636968456
transform 1 0 8372 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1636968456
transform 1 0 9476 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1636968456
transform 1 0 10580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1
transform 1 0 11684 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1636968456
transform 1 0 12420 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1636968456
transform 1 0 13524 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1636968456
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1636968456
transform 1 0 15732 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1
transform 1 0 16836 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636968456
transform 1 0 17572 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1636968456
transform 1 0 18676 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1636968456
transform 1 0 19780 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1636968456
transform 1 0 20884 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1
transform 1 0 21988 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1
transform 1 0 22540 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1636968456
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1636968456
transform 1 0 23828 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1636968456
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1636968456
transform 1 0 26036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1
transform 1 0 27140 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1
transform 1 0 27692 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1636968456
transform 1 0 27876 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1636968456
transform 1 0 28980 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1636968456
transform 1 0 30084 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1636968456
transform 1 0 31188 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1
transform 1 0 32292 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1
transform 1 0 32844 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1636968456
transform 1 0 33028 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1636968456
transform 1 0 34132 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1636968456
transform 1 0 35236 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1636968456
transform 1 0 36340 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1
transform 1 0 37444 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1
transform 1 0 37996 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1636968456
transform 1 0 38180 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1636968456
transform 1 0 39284 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1636968456
transform 1 0 40388 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1636968456
transform 1 0 41492 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1
transform 1 0 42596 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1
transform 1 0 43148 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1636968456
transform 1 0 43332 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1636968456
transform 1 0 44436 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1636968456
transform 1 0 45540 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1636968456
transform 1 0 46644 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1
transform 1 0 47748 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1
transform 1 0 48300 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1636968456
transform 1 0 48484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1636968456
transform 1 0 49588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1636968456
transform 1 0 50692 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1636968456
transform 1 0 51796 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1
transform 1 0 52900 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1
transform 1 0 53452 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1636968456
transform 1 0 53636 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1636968456
transform 1 0 54740 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1636968456
transform 1 0 55844 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1636968456
transform 1 0 56948 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1
transform 1 0 58052 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1
transform 1 0 58604 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1636968456
transform 1 0 58788 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1636968456
transform 1 0 59892 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1636968456
transform 1 0 60996 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1636968456
transform 1 0 62100 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1
transform 1 0 63204 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1
transform 1 0 63756 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1636968456
transform 1 0 63940 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1636968456
transform 1 0 65044 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1636968456
transform 1 0 66148 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1636968456
transform 1 0 67252 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1
transform 1 0 68356 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1
transform 1 0 68908 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_729
timestamp 1636968456
transform 1 0 69092 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_741
timestamp 1636968456
transform 1 0 70196 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_753
timestamp 1636968456
transform 1 0 71300 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_765
timestamp 1636968456
transform 1 0 72404 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_777
timestamp 1
transform 1 0 73508 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_783
timestamp 1
transform 1 0 74060 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_785
timestamp 1636968456
transform 1 0 74244 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_797
timestamp 1636968456
transform 1 0 75348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_809
timestamp 1636968456
transform 1 0 76452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_821
timestamp 1
transform 1 0 77556 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636968456
transform 1 0 2300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636968456
transform 1 0 3404 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636968456
transform 1 0 4692 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636968456
transform 1 0 5796 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636968456
transform 1 0 6900 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1636968456
transform 1 0 8004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1
transform 1 0 9108 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1636968456
transform 1 0 9844 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1636968456
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1636968456
transform 1 0 12052 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1636968456
transform 1 0 13156 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1
transform 1 0 14260 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636968456
transform 1 0 14996 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1636968456
transform 1 0 16100 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1636968456
transform 1 0 17204 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1636968456
transform 1 0 18308 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1
transform 1 0 19412 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1
transform 1 0 19964 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1636968456
transform 1 0 20148 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1636968456
transform 1 0 21252 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1636968456
transform 1 0 22356 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1636968456
transform 1 0 23460 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1636968456
transform 1 0 25300 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1636968456
transform 1 0 26404 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1636968456
transform 1 0 27508 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1636968456
transform 1 0 28612 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1
transform 1 0 29716 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1
transform 1 0 30268 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1636968456
transform 1 0 30452 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1636968456
transform 1 0 31556 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1636968456
transform 1 0 32660 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1636968456
transform 1 0 33764 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1
transform 1 0 34868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1
transform 1 0 35420 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1636968456
transform 1 0 35604 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1636968456
transform 1 0 36708 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1636968456
transform 1 0 37812 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1636968456
transform 1 0 38916 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1
transform 1 0 40020 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1
transform 1 0 40572 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1636968456
transform 1 0 40756 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1636968456
transform 1 0 41860 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1636968456
transform 1 0 42964 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1636968456
transform 1 0 44068 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1
transform 1 0 45172 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1
transform 1 0 45724 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1636968456
transform 1 0 45908 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1636968456
transform 1 0 47012 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1636968456
transform 1 0 48116 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1636968456
transform 1 0 49220 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1
transform 1 0 50324 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1
transform 1 0 50876 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1636968456
transform 1 0 51060 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1636968456
transform 1 0 52164 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1636968456
transform 1 0 53268 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1636968456
transform 1 0 54372 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1
transform 1 0 55476 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1
transform 1 0 56028 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1636968456
transform 1 0 56212 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1636968456
transform 1 0 57316 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1636968456
transform 1 0 58420 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1636968456
transform 1 0 59524 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1
transform 1 0 60628 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1
transform 1 0 61180 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1636968456
transform 1 0 61364 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1636968456
transform 1 0 62468 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1636968456
transform 1 0 63572 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1636968456
transform 1 0 64676 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1
transform 1 0 65780 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1
transform 1 0 66332 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1636968456
transform 1 0 66516 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1636968456
transform 1 0 67620 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_725
timestamp 1636968456
transform 1 0 68724 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_737
timestamp 1636968456
transform 1 0 69828 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_749
timestamp 1
transform 1 0 70932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_755
timestamp 1
transform 1 0 71484 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_757
timestamp 1636968456
transform 1 0 71668 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_769
timestamp 1636968456
transform 1 0 72772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_781
timestamp 1636968456
transform 1 0 73876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_793
timestamp 1636968456
transform 1 0 74980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_805
timestamp 1
transform 1 0 76084 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_811
timestamp 1
transform 1 0 76636 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_813
timestamp 1
transform 1 0 76820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_821
timestamp 1
transform 1 0 77556 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636968456
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636968456
transform 1 0 3404 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1636968456
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1636968456
transform 1 0 5612 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1
transform 1 0 6716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636968456
transform 1 0 7268 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1636968456
transform 1 0 8372 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1636968456
transform 1 0 9476 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1636968456
transform 1 0 10580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1
transform 1 0 11684 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636968456
transform 1 0 12420 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1636968456
transform 1 0 13524 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1636968456
transform 1 0 14628 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1636968456
transform 1 0 15732 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1
transform 1 0 16836 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1
transform 1 0 17388 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1636968456
transform 1 0 17572 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1636968456
transform 1 0 18676 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1636968456
transform 1 0 19780 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1636968456
transform 1 0 20884 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1
transform 1 0 21988 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1
transform 1 0 22540 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636968456
transform 1 0 22724 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636968456
transform 1 0 23828 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1636968456
transform 1 0 24932 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1636968456
transform 1 0 26036 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1
transform 1 0 27140 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1
transform 1 0 27692 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1636968456
transform 1 0 27876 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1636968456
transform 1 0 28980 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1636968456
transform 1 0 30084 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1636968456
transform 1 0 31188 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1
transform 1 0 32292 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1
transform 1 0 32844 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1636968456
transform 1 0 33028 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1636968456
transform 1 0 34132 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1636968456
transform 1 0 35236 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1636968456
transform 1 0 36340 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1
transform 1 0 37444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1
transform 1 0 37996 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1636968456
transform 1 0 38180 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1636968456
transform 1 0 39284 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1636968456
transform 1 0 40388 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1636968456
transform 1 0 41492 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1
transform 1 0 42596 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1
transform 1 0 43148 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1636968456
transform 1 0 43332 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1636968456
transform 1 0 44436 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1636968456
transform 1 0 45540 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1636968456
transform 1 0 46644 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1
transform 1 0 47748 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1
transform 1 0 48300 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1636968456
transform 1 0 48484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1636968456
transform 1 0 49588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1636968456
transform 1 0 50692 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1636968456
transform 1 0 51796 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1
transform 1 0 52900 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1
transform 1 0 53452 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1636968456
transform 1 0 53636 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1636968456
transform 1 0 54740 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1636968456
transform 1 0 55844 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1636968456
transform 1 0 56948 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1
transform 1 0 58052 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1
transform 1 0 58604 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1636968456
transform 1 0 58788 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1636968456
transform 1 0 59892 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1636968456
transform 1 0 60996 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1636968456
transform 1 0 62100 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1
transform 1 0 63204 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1
transform 1 0 63756 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1636968456
transform 1 0 63940 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1636968456
transform 1 0 65044 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1636968456
transform 1 0 66148 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1636968456
transform 1 0 67252 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1
transform 1 0 68356 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1
transform 1 0 68908 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_729
timestamp 1636968456
transform 1 0 69092 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_741
timestamp 1636968456
transform 1 0 70196 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_753
timestamp 1636968456
transform 1 0 71300 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_765
timestamp 1636968456
transform 1 0 72404 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_777
timestamp 1
transform 1 0 73508 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_783
timestamp 1
transform 1 0 74060 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_785
timestamp 1636968456
transform 1 0 74244 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_797
timestamp 1636968456
transform 1 0 75348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_809
timestamp 1636968456
transform 1 0 76452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_821
timestamp 1
transform 1 0 77556 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636968456
transform 1 0 2300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636968456
transform 1 0 3404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636968456
transform 1 0 4692 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636968456
transform 1 0 5796 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636968456
transform 1 0 6900 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1636968456
transform 1 0 8004 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1
transform 1 0 9108 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1
transform 1 0 9660 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636968456
transform 1 0 9844 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1636968456
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1636968456
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1636968456
transform 1 0 13156 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1
transform 1 0 14260 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636968456
transform 1 0 14996 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1636968456
transform 1 0 16100 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1636968456
transform 1 0 17204 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1636968456
transform 1 0 18308 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1
transform 1 0 19412 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636968456
transform 1 0 20148 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1636968456
transform 1 0 21252 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1636968456
transform 1 0 22356 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1636968456
transform 1 0 23460 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1
transform 1 0 24564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1
transform 1 0 25116 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1636968456
transform 1 0 25300 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1636968456
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1636968456
transform 1 0 27508 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1636968456
transform 1 0 28612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1
transform 1 0 29716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1
transform 1 0 30268 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1636968456
transform 1 0 30452 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1636968456
transform 1 0 31556 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1636968456
transform 1 0 32660 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1636968456
transform 1 0 33764 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1
transform 1 0 34868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1
transform 1 0 35420 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1636968456
transform 1 0 35604 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1636968456
transform 1 0 36708 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1636968456
transform 1 0 37812 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1636968456
transform 1 0 38916 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1
transform 1 0 40020 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1
transform 1 0 40572 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1636968456
transform 1 0 40756 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1636968456
transform 1 0 41860 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1636968456
transform 1 0 42964 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1636968456
transform 1 0 44068 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1
transform 1 0 45172 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1
transform 1 0 45724 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1636968456
transform 1 0 45908 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1636968456
transform 1 0 47012 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1636968456
transform 1 0 48116 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1636968456
transform 1 0 49220 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1
transform 1 0 50324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1
transform 1 0 50876 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1636968456
transform 1 0 51060 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1636968456
transform 1 0 52164 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1636968456
transform 1 0 53268 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1636968456
transform 1 0 54372 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1
transform 1 0 55476 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1
transform 1 0 56028 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1636968456
transform 1 0 56212 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1636968456
transform 1 0 57316 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1636968456
transform 1 0 58420 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1636968456
transform 1 0 59524 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1
transform 1 0 60628 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1
transform 1 0 61180 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1636968456
transform 1 0 61364 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1636968456
transform 1 0 62468 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1636968456
transform 1 0 63572 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1636968456
transform 1 0 64676 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1
transform 1 0 65780 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1
transform 1 0 66332 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1636968456
transform 1 0 66516 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1636968456
transform 1 0 67620 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_725
timestamp 1636968456
transform 1 0 68724 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_737
timestamp 1636968456
transform 1 0 69828 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_749
timestamp 1
transform 1 0 70932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 1
transform 1 0 71484 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_757
timestamp 1636968456
transform 1 0 71668 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_769
timestamp 1636968456
transform 1 0 72772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_781
timestamp 1636968456
transform 1 0 73876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_793
timestamp 1636968456
transform 1 0 74980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_805
timestamp 1
transform 1 0 76084 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_811
timestamp 1
transform 1 0 76636 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_813
timestamp 1
transform 1 0 76820 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636968456
transform 1 0 2300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636968456
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636968456
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636968456
transform 1 0 5612 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1
transform 1 0 6716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1
transform 1 0 7084 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636968456
transform 1 0 7268 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1636968456
transform 1 0 8372 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1636968456
transform 1 0 9476 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1636968456
transform 1 0 10580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1
transform 1 0 11684 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1636968456
transform 1 0 12420 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1636968456
transform 1 0 13524 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1636968456
transform 1 0 14628 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1636968456
transform 1 0 15732 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1
transform 1 0 16836 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1
transform 1 0 17388 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1636968456
transform 1 0 17572 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1636968456
transform 1 0 18676 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1636968456
transform 1 0 19780 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1636968456
transform 1 0 20884 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1
transform 1 0 21988 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1
transform 1 0 22540 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1636968456
transform 1 0 22724 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1636968456
transform 1 0 23828 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1636968456
transform 1 0 24932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1636968456
transform 1 0 26036 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1
transform 1 0 27140 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1
transform 1 0 27692 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1636968456
transform 1 0 27876 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1636968456
transform 1 0 28980 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1636968456
transform 1 0 30084 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1636968456
transform 1 0 31188 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1
transform 1 0 32292 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1
transform 1 0 32844 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1636968456
transform 1 0 33028 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1636968456
transform 1 0 34132 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1636968456
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1636968456
transform 1 0 36340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1
transform 1 0 37444 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1
transform 1 0 37996 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1636968456
transform 1 0 38180 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1636968456
transform 1 0 39284 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1636968456
transform 1 0 40388 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1636968456
transform 1 0 41492 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1
transform 1 0 42596 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1
transform 1 0 43148 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1636968456
transform 1 0 43332 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1636968456
transform 1 0 44436 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1636968456
transform 1 0 45540 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1636968456
transform 1 0 46644 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1
transform 1 0 47748 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1
transform 1 0 48300 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1636968456
transform 1 0 48484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1636968456
transform 1 0 49588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1636968456
transform 1 0 50692 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1636968456
transform 1 0 51796 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1
transform 1 0 52900 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1
transform 1 0 53452 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1636968456
transform 1 0 53636 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1636968456
transform 1 0 54740 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1636968456
transform 1 0 55844 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1636968456
transform 1 0 56948 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1
transform 1 0 58052 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1
transform 1 0 58604 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1636968456
transform 1 0 58788 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1636968456
transform 1 0 59892 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1636968456
transform 1 0 60996 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1636968456
transform 1 0 62100 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1
transform 1 0 63204 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1
transform 1 0 63756 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1636968456
transform 1 0 63940 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1636968456
transform 1 0 65044 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1636968456
transform 1 0 66148 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1636968456
transform 1 0 67252 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1
transform 1 0 68356 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1
transform 1 0 68908 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_729
timestamp 1636968456
transform 1 0 69092 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_741
timestamp 1636968456
transform 1 0 70196 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_753
timestamp 1636968456
transform 1 0 71300 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_765
timestamp 1636968456
transform 1 0 72404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_777
timestamp 1
transform 1 0 73508 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_783
timestamp 1
transform 1 0 74060 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_785
timestamp 1636968456
transform 1 0 74244 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_797
timestamp 1636968456
transform 1 0 75348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_809
timestamp 1636968456
transform 1 0 76452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_821
timestamp 1
transform 1 0 77556 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636968456
transform 1 0 2300 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636968456
transform 1 0 3404 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636968456
transform 1 0 4692 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636968456
transform 1 0 5796 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636968456
transform 1 0 6900 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1636968456
transform 1 0 8004 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1
transform 1 0 9108 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1636968456
transform 1 0 9844 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1636968456
transform 1 0 10948 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1636968456
transform 1 0 12052 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1636968456
transform 1 0 13156 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1
transform 1 0 14260 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1
transform 1 0 14812 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1636968456
transform 1 0 14996 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1636968456
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1636968456
transform 1 0 17204 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1636968456
transform 1 0 18308 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1
transform 1 0 19412 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1636968456
transform 1 0 20148 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1636968456
transform 1 0 21252 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1636968456
transform 1 0 22356 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1636968456
transform 1 0 23460 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1
transform 1 0 24564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1
transform 1 0 25116 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1636968456
transform 1 0 25300 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1636968456
transform 1 0 26404 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1636968456
transform 1 0 27508 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1636968456
transform 1 0 28612 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1
transform 1 0 29716 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1
transform 1 0 30268 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1636968456
transform 1 0 30452 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1636968456
transform 1 0 31556 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1636968456
transform 1 0 32660 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1636968456
transform 1 0 33764 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1
transform 1 0 34868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1
transform 1 0 35420 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1636968456
transform 1 0 35604 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1636968456
transform 1 0 36708 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1636968456
transform 1 0 37812 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1636968456
transform 1 0 38916 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1
transform 1 0 40020 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1
transform 1 0 40572 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1636968456
transform 1 0 40756 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1636968456
transform 1 0 41860 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1636968456
transform 1 0 42964 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1636968456
transform 1 0 44068 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1
transform 1 0 45172 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1
transform 1 0 45724 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1636968456
transform 1 0 45908 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1636968456
transform 1 0 47012 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1636968456
transform 1 0 48116 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1636968456
transform 1 0 49220 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1
transform 1 0 50324 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1
transform 1 0 50876 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1636968456
transform 1 0 51060 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1636968456
transform 1 0 52164 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1636968456
transform 1 0 53268 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1636968456
transform 1 0 54372 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1
transform 1 0 55476 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1
transform 1 0 56028 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1636968456
transform 1 0 56212 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1636968456
transform 1 0 57316 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1636968456
transform 1 0 58420 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1636968456
transform 1 0 59524 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1
transform 1 0 60628 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1
transform 1 0 61180 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1636968456
transform 1 0 61364 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1636968456
transform 1 0 62468 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1636968456
transform 1 0 63572 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1636968456
transform 1 0 64676 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1
transform 1 0 65780 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1
transform 1 0 66332 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1636968456
transform 1 0 66516 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1636968456
transform 1 0 67620 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_725
timestamp 1636968456
transform 1 0 68724 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_737
timestamp 1636968456
transform 1 0 69828 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_749
timestamp 1
transform 1 0 70932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_755
timestamp 1
transform 1 0 71484 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_757
timestamp 1636968456
transform 1 0 71668 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_769
timestamp 1636968456
transform 1 0 72772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_781
timestamp 1636968456
transform 1 0 73876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_793
timestamp 1636968456
transform 1 0 74980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_805
timestamp 1
transform 1 0 76084 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_811
timestamp 1
transform 1 0 76636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_813
timestamp 1
transform 1 0 76820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_821
timestamp 1
transform 1 0 77556 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636968456
transform 1 0 2300 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636968456
transform 1 0 3404 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636968456
transform 1 0 4508 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636968456
transform 1 0 5612 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1
transform 1 0 6716 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1
transform 1 0 7084 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636968456
transform 1 0 7268 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1636968456
transform 1 0 8372 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1636968456
transform 1 0 9476 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1636968456
transform 1 0 10580 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1
transform 1 0 11684 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1
transform 1 0 12236 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1636968456
transform 1 0 12420 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1636968456
transform 1 0 13524 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1636968456
transform 1 0 14628 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1636968456
transform 1 0 15732 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1
transform 1 0 16836 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1
transform 1 0 17388 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1636968456
transform 1 0 17572 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1636968456
transform 1 0 18676 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1636968456
transform 1 0 19780 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1636968456
transform 1 0 20884 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1
transform 1 0 21988 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1
transform 1 0 22540 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1636968456
transform 1 0 22724 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1636968456
transform 1 0 23828 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1636968456
transform 1 0 24932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1636968456
transform 1 0 26036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1
transform 1 0 27140 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1
transform 1 0 27692 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1636968456
transform 1 0 27876 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1636968456
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1636968456
transform 1 0 30084 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1636968456
transform 1 0 31188 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1
transform 1 0 32292 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1
transform 1 0 32844 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1636968456
transform 1 0 33028 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1636968456
transform 1 0 34132 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1636968456
transform 1 0 35236 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1636968456
transform 1 0 36340 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1
transform 1 0 37444 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1
transform 1 0 37996 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1636968456
transform 1 0 38180 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1636968456
transform 1 0 39284 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1636968456
transform 1 0 40388 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1636968456
transform 1 0 41492 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1
transform 1 0 42596 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1
transform 1 0 43148 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1636968456
transform 1 0 43332 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1636968456
transform 1 0 44436 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1636968456
transform 1 0 45540 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1636968456
transform 1 0 46644 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1
transform 1 0 47748 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1
transform 1 0 48300 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1636968456
transform 1 0 48484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1636968456
transform 1 0 49588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1636968456
transform 1 0 50692 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1636968456
transform 1 0 51796 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1
transform 1 0 52900 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1
transform 1 0 53452 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1636968456
transform 1 0 53636 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1636968456
transform 1 0 54740 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1636968456
transform 1 0 55844 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1636968456
transform 1 0 56948 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1
transform 1 0 58052 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1
transform 1 0 58604 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1636968456
transform 1 0 58788 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1636968456
transform 1 0 59892 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1636968456
transform 1 0 60996 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1636968456
transform 1 0 62100 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1
transform 1 0 63204 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1
transform 1 0 63756 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1636968456
transform 1 0 63940 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1636968456
transform 1 0 65044 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1636968456
transform 1 0 66148 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1636968456
transform 1 0 67252 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1
transform 1 0 68356 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1
transform 1 0 68908 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_729
timestamp 1636968456
transform 1 0 69092 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_741
timestamp 1636968456
transform 1 0 70196 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_753
timestamp 1636968456
transform 1 0 71300 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_765
timestamp 1636968456
transform 1 0 72404 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_777
timestamp 1
transform 1 0 73508 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 1
transform 1 0 74060 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_785
timestamp 1636968456
transform 1 0 74244 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_797
timestamp 1636968456
transform 1 0 75348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_809
timestamp 1636968456
transform 1 0 76452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_821
timestamp 1
transform 1 0 77556 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636968456
transform 1 0 3404 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 4508 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636968456
transform 1 0 4692 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636968456
transform 1 0 5796 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636968456
transform 1 0 6900 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1636968456
transform 1 0 8004 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1
transform 1 0 9108 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1
transform 1 0 9660 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1636968456
transform 1 0 9844 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1636968456
transform 1 0 10948 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1636968456
transform 1 0 12052 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1636968456
transform 1 0 13156 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1
transform 1 0 14260 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1
transform 1 0 14812 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1636968456
transform 1 0 14996 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1636968456
transform 1 0 16100 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1636968456
transform 1 0 17204 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1636968456
transform 1 0 18308 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1
transform 1 0 19412 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1
transform 1 0 19964 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1636968456
transform 1 0 20148 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1636968456
transform 1 0 21252 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1636968456
transform 1 0 22356 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1636968456
transform 1 0 23460 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1
transform 1 0 24564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1
transform 1 0 25116 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636968456
transform 1 0 25300 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1636968456
transform 1 0 26404 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1636968456
transform 1 0 27508 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1636968456
transform 1 0 28612 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1
transform 1 0 29716 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1
transform 1 0 30268 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1636968456
transform 1 0 30452 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1636968456
transform 1 0 31556 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1636968456
transform 1 0 32660 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1636968456
transform 1 0 33764 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1
transform 1 0 34868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1
transform 1 0 35420 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1636968456
transform 1 0 35604 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1636968456
transform 1 0 36708 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1636968456
transform 1 0 37812 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1636968456
transform 1 0 38916 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1
transform 1 0 40020 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1
transform 1 0 40572 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1636968456
transform 1 0 40756 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1636968456
transform 1 0 41860 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1636968456
transform 1 0 42964 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1636968456
transform 1 0 44068 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1
transform 1 0 45172 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1
transform 1 0 45724 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1636968456
transform 1 0 45908 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1636968456
transform 1 0 47012 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1636968456
transform 1 0 48116 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1636968456
transform 1 0 49220 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1
transform 1 0 50324 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1
transform 1 0 50876 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1636968456
transform 1 0 51060 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1636968456
transform 1 0 52164 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1636968456
transform 1 0 53268 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1636968456
transform 1 0 54372 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1
transform 1 0 55476 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1
transform 1 0 56028 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1636968456
transform 1 0 56212 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1636968456
transform 1 0 57316 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1636968456
transform 1 0 58420 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1636968456
transform 1 0 59524 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1
transform 1 0 60628 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1
transform 1 0 61180 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1636968456
transform 1 0 61364 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1636968456
transform 1 0 62468 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1636968456
transform 1 0 63572 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1636968456
transform 1 0 64676 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1
transform 1 0 65780 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1
transform 1 0 66332 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1636968456
transform 1 0 66516 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1636968456
transform 1 0 67620 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_725
timestamp 1636968456
transform 1 0 68724 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_737
timestamp 1636968456
transform 1 0 69828 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 1
transform 1 0 70932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 1
transform 1 0 71484 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_757
timestamp 1636968456
transform 1 0 71668 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_769
timestamp 1636968456
transform 1 0 72772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_781
timestamp 1636968456
transform 1 0 73876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_793
timestamp 1636968456
transform 1 0 74980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 1
transform 1 0 76084 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 1
transform 1 0 76636 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_813
timestamp 1
transform 1 0 76820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_821
timestamp 1
transform 1 0 77556 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636968456
transform 1 0 2300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636968456
transform 1 0 3404 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636968456
transform 1 0 4508 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636968456
transform 1 0 5612 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1
transform 1 0 6716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1
transform 1 0 7084 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636968456
transform 1 0 7268 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1636968456
transform 1 0 8372 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1636968456
transform 1 0 9476 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1636968456
transform 1 0 10580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1
transform 1 0 11684 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1636968456
transform 1 0 12420 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1636968456
transform 1 0 13524 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1636968456
transform 1 0 14628 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1636968456
transform 1 0 15732 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1
transform 1 0 16836 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1
transform 1 0 17388 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1636968456
transform 1 0 17572 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1636968456
transform 1 0 18676 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1636968456
transform 1 0 19780 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1636968456
transform 1 0 20884 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1
transform 1 0 21988 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1
transform 1 0 22540 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636968456
transform 1 0 22724 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1636968456
transform 1 0 23828 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1636968456
transform 1 0 24932 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1636968456
transform 1 0 26036 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1
transform 1 0 27140 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1
transform 1 0 27692 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1636968456
transform 1 0 27876 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1636968456
transform 1 0 28980 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1636968456
transform 1 0 30084 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1636968456
transform 1 0 31188 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1
transform 1 0 32292 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1
transform 1 0 32844 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1636968456
transform 1 0 33028 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1636968456
transform 1 0 34132 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1636968456
transform 1 0 35236 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1636968456
transform 1 0 36340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1
transform 1 0 37444 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1
transform 1 0 37996 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1636968456
transform 1 0 38180 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1636968456
transform 1 0 39284 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1636968456
transform 1 0 40388 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1636968456
transform 1 0 41492 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1
transform 1 0 42596 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1
transform 1 0 43148 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1636968456
transform 1 0 43332 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1636968456
transform 1 0 44436 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1636968456
transform 1 0 45540 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1636968456
transform 1 0 46644 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1
transform 1 0 47748 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1
transform 1 0 48300 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1636968456
transform 1 0 48484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1636968456
transform 1 0 49588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1636968456
transform 1 0 50692 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1636968456
transform 1 0 51796 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1
transform 1 0 52900 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1
transform 1 0 53452 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1636968456
transform 1 0 53636 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1636968456
transform 1 0 54740 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1636968456
transform 1 0 55844 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1636968456
transform 1 0 56948 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1
transform 1 0 58052 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1
transform 1 0 58604 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1636968456
transform 1 0 58788 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1636968456
transform 1 0 59892 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1636968456
transform 1 0 60996 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1636968456
transform 1 0 62100 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1
transform 1 0 63204 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1
transform 1 0 63756 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1636968456
transform 1 0 63940 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1636968456
transform 1 0 65044 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1636968456
transform 1 0 66148 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1636968456
transform 1 0 67252 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1
transform 1 0 68356 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1
transform 1 0 68908 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_729
timestamp 1636968456
transform 1 0 69092 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_741
timestamp 1636968456
transform 1 0 70196 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_753
timestamp 1636968456
transform 1 0 71300 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_765
timestamp 1636968456
transform 1 0 72404 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_777
timestamp 1
transform 1 0 73508 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 1
transform 1 0 74060 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_785
timestamp 1636968456
transform 1 0 74244 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_797
timestamp 1636968456
transform 1 0 75348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_809
timestamp 1636968456
transform 1 0 76452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_821
timestamp 1
transform 1 0 77556 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636968456
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636968456
transform 1 0 3404 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636968456
transform 1 0 4692 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636968456
transform 1 0 5796 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636968456
transform 1 0 6900 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1636968456
transform 1 0 8004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1
transform 1 0 9108 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1
transform 1 0 9660 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1636968456
transform 1 0 9844 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1636968456
transform 1 0 10948 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1636968456
transform 1 0 12052 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1636968456
transform 1 0 13156 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1
transform 1 0 14260 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1
transform 1 0 14812 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1636968456
transform 1 0 14996 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1636968456
transform 1 0 16100 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1636968456
transform 1 0 17204 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1636968456
transform 1 0 18308 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1
transform 1 0 19412 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1
transform 1 0 19964 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1636968456
transform 1 0 20148 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1636968456
transform 1 0 21252 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1636968456
transform 1 0 22356 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1636968456
transform 1 0 23460 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1
transform 1 0 24564 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1
transform 1 0 25116 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636968456
transform 1 0 25300 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1636968456
transform 1 0 26404 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1636968456
transform 1 0 27508 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1636968456
transform 1 0 28612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1
transform 1 0 29716 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1
transform 1 0 30268 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1636968456
transform 1 0 30452 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1636968456
transform 1 0 31556 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1636968456
transform 1 0 32660 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1636968456
transform 1 0 33764 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1
transform 1 0 34868 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1
transform 1 0 35420 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1636968456
transform 1 0 35604 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1636968456
transform 1 0 36708 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1636968456
transform 1 0 37812 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1636968456
transform 1 0 38916 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1
transform 1 0 40020 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1
transform 1 0 40572 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1636968456
transform 1 0 40756 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1636968456
transform 1 0 41860 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1636968456
transform 1 0 42964 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1636968456
transform 1 0 44068 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1
transform 1 0 45172 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1
transform 1 0 45724 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1636968456
transform 1 0 45908 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1636968456
transform 1 0 47012 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1636968456
transform 1 0 48116 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1636968456
transform 1 0 49220 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1
transform 1 0 50324 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1
transform 1 0 50876 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1636968456
transform 1 0 51060 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1636968456
transform 1 0 52164 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1636968456
transform 1 0 53268 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1636968456
transform 1 0 54372 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1
transform 1 0 55476 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1
transform 1 0 56028 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1636968456
transform 1 0 56212 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1636968456
transform 1 0 57316 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1636968456
transform 1 0 58420 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1636968456
transform 1 0 59524 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1
transform 1 0 60628 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1
transform 1 0 61180 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1636968456
transform 1 0 61364 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1636968456
transform 1 0 62468 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1636968456
transform 1 0 63572 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1636968456
transform 1 0 64676 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1
transform 1 0 65780 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1
transform 1 0 66332 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1636968456
transform 1 0 66516 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1636968456
transform 1 0 67620 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_725
timestamp 1636968456
transform 1 0 68724 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_737
timestamp 1636968456
transform 1 0 69828 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_749
timestamp 1
transform 1 0 70932 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 1
transform 1 0 71484 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_757
timestamp 1636968456
transform 1 0 71668 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_769
timestamp 1636968456
transform 1 0 72772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_781
timestamp 1636968456
transform 1 0 73876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_793
timestamp 1636968456
transform 1 0 74980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_805
timestamp 1
transform 1 0 76084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 1
transform 1 0 76636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_813
timestamp 1
transform 1 0 76820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_821
timestamp 1
transform 1 0 77556 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636968456
transform 1 0 2300 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636968456
transform 1 0 3404 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1636968456
transform 1 0 4508 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1636968456
transform 1 0 5612 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1
transform 1 0 6716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1
transform 1 0 7084 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636968456
transform 1 0 7268 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1636968456
transform 1 0 8372 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1636968456
transform 1 0 9476 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1636968456
transform 1 0 10580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1
transform 1 0 11684 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1636968456
transform 1 0 12420 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1636968456
transform 1 0 13524 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1636968456
transform 1 0 14628 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1636968456
transform 1 0 15732 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1
transform 1 0 16836 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1
transform 1 0 17388 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1636968456
transform 1 0 17572 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1636968456
transform 1 0 18676 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1636968456
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1636968456
transform 1 0 20884 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1
transform 1 0 21988 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1
transform 1 0 22540 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1636968456
transform 1 0 22724 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1636968456
transform 1 0 23828 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1636968456
transform 1 0 24932 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1636968456
transform 1 0 26036 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1
transform 1 0 27140 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1
transform 1 0 27692 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1636968456
transform 1 0 27876 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1636968456
transform 1 0 28980 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1636968456
transform 1 0 30084 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1636968456
transform 1 0 31188 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1
transform 1 0 32292 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1
transform 1 0 32844 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1636968456
transform 1 0 33028 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1636968456
transform 1 0 34132 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1636968456
transform 1 0 35236 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1636968456
transform 1 0 36340 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1
transform 1 0 37444 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1
transform 1 0 37996 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1636968456
transform 1 0 38180 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1636968456
transform 1 0 39284 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1636968456
transform 1 0 40388 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1636968456
transform 1 0 41492 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1
transform 1 0 42596 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1
transform 1 0 43148 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1636968456
transform 1 0 43332 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1636968456
transform 1 0 44436 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1636968456
transform 1 0 45540 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1636968456
transform 1 0 46644 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1
transform 1 0 47748 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1
transform 1 0 48300 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1636968456
transform 1 0 48484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1636968456
transform 1 0 49588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1636968456
transform 1 0 50692 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1636968456
transform 1 0 51796 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1
transform 1 0 52900 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1
transform 1 0 53452 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1636968456
transform 1 0 53636 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1636968456
transform 1 0 54740 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1636968456
transform 1 0 55844 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1636968456
transform 1 0 56948 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1
transform 1 0 58052 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1
transform 1 0 58604 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1636968456
transform 1 0 58788 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1636968456
transform 1 0 59892 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1636968456
transform 1 0 60996 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1636968456
transform 1 0 62100 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1
transform 1 0 63204 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1
transform 1 0 63756 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1636968456
transform 1 0 63940 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1636968456
transform 1 0 65044 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1636968456
transform 1 0 66148 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1636968456
transform 1 0 67252 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1
transform 1 0 68356 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1
transform 1 0 68908 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_729
timestamp 1636968456
transform 1 0 69092 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_741
timestamp 1636968456
transform 1 0 70196 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_753
timestamp 1636968456
transform 1 0 71300 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_765
timestamp 1636968456
transform 1 0 72404 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_777
timestamp 1
transform 1 0 73508 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_783
timestamp 1
transform 1 0 74060 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_785
timestamp 1636968456
transform 1 0 74244 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_797
timestamp 1636968456
transform 1 0 75348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_809
timestamp 1636968456
transform 1 0 76452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_821
timestamp 1
transform 1 0 77556 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636968456
transform 1 0 2300 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636968456
transform 1 0 3404 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1636968456
transform 1 0 4692 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1636968456
transform 1 0 5796 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1636968456
transform 1 0 6900 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1636968456
transform 1 0 8004 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1
transform 1 0 9108 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1636968456
transform 1 0 9844 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1636968456
transform 1 0 10948 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1636968456
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1636968456
transform 1 0 13156 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1
transform 1 0 14260 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1
transform 1 0 14812 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1636968456
transform 1 0 14996 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1636968456
transform 1 0 16100 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1636968456
transform 1 0 17204 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1636968456
transform 1 0 18308 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1
transform 1 0 19412 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1
transform 1 0 19964 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1636968456
transform 1 0 20148 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1636968456
transform 1 0 21252 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1636968456
transform 1 0 22356 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1636968456
transform 1 0 23460 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1
transform 1 0 24564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1
transform 1 0 25116 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1636968456
transform 1 0 25300 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1636968456
transform 1 0 26404 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1636968456
transform 1 0 27508 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1636968456
transform 1 0 28612 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1
transform 1 0 29716 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1
transform 1 0 30268 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1636968456
transform 1 0 30452 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1636968456
transform 1 0 31556 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1636968456
transform 1 0 32660 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1636968456
transform 1 0 33764 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1
transform 1 0 34868 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1
transform 1 0 35420 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1636968456
transform 1 0 35604 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1636968456
transform 1 0 36708 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1636968456
transform 1 0 37812 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1636968456
transform 1 0 38916 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1
transform 1 0 40020 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1
transform 1 0 40572 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1636968456
transform 1 0 40756 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1636968456
transform 1 0 41860 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1636968456
transform 1 0 42964 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1636968456
transform 1 0 44068 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1
transform 1 0 45172 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1
transform 1 0 45724 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1636968456
transform 1 0 45908 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1636968456
transform 1 0 47012 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1636968456
transform 1 0 48116 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1636968456
transform 1 0 49220 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1
transform 1 0 50324 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1
transform 1 0 50876 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1636968456
transform 1 0 51060 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1636968456
transform 1 0 52164 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1636968456
transform 1 0 53268 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1636968456
transform 1 0 54372 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1
transform 1 0 55476 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1
transform 1 0 56028 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1636968456
transform 1 0 56212 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1636968456
transform 1 0 57316 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1636968456
transform 1 0 58420 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1636968456
transform 1 0 59524 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1
transform 1 0 60628 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1
transform 1 0 61180 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1636968456
transform 1 0 61364 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1636968456
transform 1 0 62468 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1636968456
transform 1 0 63572 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1636968456
transform 1 0 64676 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1
transform 1 0 65780 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1
transform 1 0 66332 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1636968456
transform 1 0 66516 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1636968456
transform 1 0 67620 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_725
timestamp 1636968456
transform 1 0 68724 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_737
timestamp 1636968456
transform 1 0 69828 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 1
transform 1 0 70932 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 1
transform 1 0 71484 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_757
timestamp 1636968456
transform 1 0 71668 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_769
timestamp 1636968456
transform 1 0 72772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_781
timestamp 1636968456
transform 1 0 73876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_793
timestamp 1636968456
transform 1 0 74980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_805
timestamp 1
transform 1 0 76084 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 1
transform 1 0 76636 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_813
timestamp 1
transform 1 0 76820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_821
timestamp 1
transform 1 0 77556 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636968456
transform 1 0 2300 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636968456
transform 1 0 3404 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1636968456
transform 1 0 4508 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1636968456
transform 1 0 5612 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1
transform 1 0 6716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1
transform 1 0 7084 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636968456
transform 1 0 7268 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1636968456
transform 1 0 8372 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1636968456
transform 1 0 9476 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1636968456
transform 1 0 10580 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1
transform 1 0 11684 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1
transform 1 0 12236 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1636968456
transform 1 0 12420 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1636968456
transform 1 0 13524 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1636968456
transform 1 0 14628 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1636968456
transform 1 0 15732 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1
transform 1 0 16836 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1
transform 1 0 17388 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1636968456
transform 1 0 17572 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1636968456
transform 1 0 18676 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1636968456
transform 1 0 19780 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1636968456
transform 1 0 20884 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1
transform 1 0 21988 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1
transform 1 0 22540 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1636968456
transform 1 0 22724 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1636968456
transform 1 0 23828 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1636968456
transform 1 0 24932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1636968456
transform 1 0 26036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1
transform 1 0 27140 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1
transform 1 0 27692 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1636968456
transform 1 0 27876 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1636968456
transform 1 0 28980 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1636968456
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1636968456
transform 1 0 31188 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1
transform 1 0 32292 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1
transform 1 0 32844 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1636968456
transform 1 0 33028 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1636968456
transform 1 0 34132 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1636968456
transform 1 0 35236 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1636968456
transform 1 0 36340 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1
transform 1 0 37444 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1
transform 1 0 37996 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1636968456
transform 1 0 38180 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1636968456
transform 1 0 39284 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1636968456
transform 1 0 40388 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1636968456
transform 1 0 41492 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1
transform 1 0 42596 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1
transform 1 0 43148 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1636968456
transform 1 0 43332 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1636968456
transform 1 0 44436 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1636968456
transform 1 0 45540 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1636968456
transform 1 0 46644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1
transform 1 0 47748 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1
transform 1 0 48300 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1636968456
transform 1 0 48484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1636968456
transform 1 0 49588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1636968456
transform 1 0 50692 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1636968456
transform 1 0 51796 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1
transform 1 0 52900 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1
transform 1 0 53452 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1636968456
transform 1 0 53636 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1636968456
transform 1 0 54740 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1636968456
transform 1 0 55844 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1636968456
transform 1 0 56948 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1
transform 1 0 58052 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1
transform 1 0 58604 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1636968456
transform 1 0 58788 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1636968456
transform 1 0 59892 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1636968456
transform 1 0 60996 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1636968456
transform 1 0 62100 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1
transform 1 0 63204 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1
transform 1 0 63756 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1636968456
transform 1 0 63940 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1636968456
transform 1 0 65044 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1636968456
transform 1 0 66148 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1636968456
transform 1 0 67252 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1
transform 1 0 68356 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1
transform 1 0 68908 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_729
timestamp 1636968456
transform 1 0 69092 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_741
timestamp 1636968456
transform 1 0 70196 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_753
timestamp 1636968456
transform 1 0 71300 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_765
timestamp 1636968456
transform 1 0 72404 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_777
timestamp 1
transform 1 0 73508 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_783
timestamp 1
transform 1 0 74060 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_785
timestamp 1636968456
transform 1 0 74244 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_797
timestamp 1636968456
transform 1 0 75348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_809
timestamp 1
transform 1 0 76452 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_817
timestamp 1
transform 1 0 77188 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636968456
transform 1 0 2300 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636968456
transform 1 0 3404 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 4508 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636968456
transform 1 0 4692 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1636968456
transform 1 0 5796 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1636968456
transform 1 0 6900 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1636968456
transform 1 0 8004 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1
transform 1 0 9108 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1
transform 1 0 9660 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1636968456
transform 1 0 9844 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1636968456
transform 1 0 10948 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1636968456
transform 1 0 12052 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1636968456
transform 1 0 13156 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1
transform 1 0 14260 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1
transform 1 0 14812 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1636968456
transform 1 0 14996 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1636968456
transform 1 0 16100 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1636968456
transform 1 0 17204 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1636968456
transform 1 0 18308 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1
transform 1 0 19412 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1
transform 1 0 19964 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1636968456
transform 1 0 20148 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1636968456
transform 1 0 21252 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1636968456
transform 1 0 22356 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1636968456
transform 1 0 23460 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1
transform 1 0 24564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1
transform 1 0 25116 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1636968456
transform 1 0 25300 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1636968456
transform 1 0 26404 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1636968456
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1636968456
transform 1 0 28612 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1
transform 1 0 29716 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1
transform 1 0 30268 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1636968456
transform 1 0 30452 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1636968456
transform 1 0 31556 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1636968456
transform 1 0 32660 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1636968456
transform 1 0 33764 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1
transform 1 0 34868 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1
transform 1 0 35420 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1636968456
transform 1 0 35604 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1636968456
transform 1 0 36708 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1636968456
transform 1 0 37812 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1636968456
transform 1 0 38916 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1
transform 1 0 40020 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1
transform 1 0 40572 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1636968456
transform 1 0 40756 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1636968456
transform 1 0 41860 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1636968456
transform 1 0 42964 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1636968456
transform 1 0 44068 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1
transform 1 0 45172 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1
transform 1 0 45724 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1636968456
transform 1 0 45908 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1636968456
transform 1 0 47012 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1636968456
transform 1 0 48116 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1636968456
transform 1 0 49220 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1
transform 1 0 50324 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1
transform 1 0 50876 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1636968456
transform 1 0 51060 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1636968456
transform 1 0 52164 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1636968456
transform 1 0 53268 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1636968456
transform 1 0 54372 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1
transform 1 0 55476 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1
transform 1 0 56028 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1636968456
transform 1 0 56212 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1636968456
transform 1 0 57316 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1636968456
transform 1 0 58420 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1636968456
transform 1 0 59524 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1
transform 1 0 60628 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1
transform 1 0 61180 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1636968456
transform 1 0 61364 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1636968456
transform 1 0 62468 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1636968456
transform 1 0 63572 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1636968456
transform 1 0 64676 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1
transform 1 0 65780 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1
transform 1 0 66332 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1636968456
transform 1 0 66516 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1636968456
transform 1 0 67620 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_725
timestamp 1636968456
transform 1 0 68724 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_737
timestamp 1636968456
transform 1 0 69828 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_749
timestamp 1
transform 1 0 70932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_755
timestamp 1
transform 1 0 71484 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_757
timestamp 1636968456
transform 1 0 71668 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_769
timestamp 1636968456
transform 1 0 72772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_781
timestamp 1636968456
transform 1 0 73876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_793
timestamp 1636968456
transform 1 0 74980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 1
transform 1 0 76084 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 1
transform 1 0 76636 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_813
timestamp 1
transform 1 0 76820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_821
timestamp 1
transform 1 0 77556 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1636968456
transform 1 0 2300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1636968456
transform 1 0 3404 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1636968456
transform 1 0 4508 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1636968456
transform 1 0 5612 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1
transform 1 0 6716 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1
transform 1 0 7084 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636968456
transform 1 0 7268 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1636968456
transform 1 0 8372 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1636968456
transform 1 0 9476 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1636968456
transform 1 0 10580 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1
transform 1 0 11684 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1
transform 1 0 12236 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1636968456
transform 1 0 12420 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1636968456
transform 1 0 13524 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1636968456
transform 1 0 14628 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1636968456
transform 1 0 15732 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1
transform 1 0 16836 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1
transform 1 0 17388 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1636968456
transform 1 0 17572 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1636968456
transform 1 0 18676 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1636968456
transform 1 0 19780 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1636968456
transform 1 0 20884 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1
transform 1 0 21988 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1
transform 1 0 22540 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1636968456
transform 1 0 22724 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1636968456
transform 1 0 23828 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1636968456
transform 1 0 24932 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1636968456
transform 1 0 26036 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1
transform 1 0 27140 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1
transform 1 0 27692 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1636968456
transform 1 0 27876 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1636968456
transform 1 0 28980 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1636968456
transform 1 0 30084 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1636968456
transform 1 0 31188 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1
transform 1 0 32292 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1
transform 1 0 32844 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1636968456
transform 1 0 33028 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1636968456
transform 1 0 34132 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1636968456
transform 1 0 35236 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1636968456
transform 1 0 36340 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1
transform 1 0 37444 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1
transform 1 0 37996 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1636968456
transform 1 0 38180 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1636968456
transform 1 0 39284 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1636968456
transform 1 0 40388 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1636968456
transform 1 0 41492 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1
transform 1 0 42596 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1
transform 1 0 43148 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1636968456
transform 1 0 43332 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1636968456
transform 1 0 44436 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1636968456
transform 1 0 45540 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1636968456
transform 1 0 46644 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1
transform 1 0 47748 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1
transform 1 0 48300 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1636968456
transform 1 0 48484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1636968456
transform 1 0 49588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1636968456
transform 1 0 50692 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1636968456
transform 1 0 51796 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1
transform 1 0 52900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1
transform 1 0 53452 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1636968456
transform 1 0 53636 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1636968456
transform 1 0 54740 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1636968456
transform 1 0 55844 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1636968456
transform 1 0 56948 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1
transform 1 0 58052 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1
transform 1 0 58604 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1636968456
transform 1 0 58788 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1636968456
transform 1 0 59892 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1636968456
transform 1 0 60996 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1636968456
transform 1 0 62100 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1
transform 1 0 63204 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1
transform 1 0 63756 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1636968456
transform 1 0 63940 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1636968456
transform 1 0 65044 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1636968456
transform 1 0 66148 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1636968456
transform 1 0 67252 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1
transform 1 0 68356 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1
transform 1 0 68908 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_729
timestamp 1636968456
transform 1 0 69092 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_741
timestamp 1636968456
transform 1 0 70196 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_753
timestamp 1636968456
transform 1 0 71300 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_765
timestamp 1636968456
transform 1 0 72404 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 1
transform 1 0 73508 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 1
transform 1 0 74060 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_785
timestamp 1636968456
transform 1 0 74244 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_797
timestamp 1636968456
transform 1 0 75348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_809
timestamp 1636968456
transform 1 0 76452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_821
timestamp 1
transform 1 0 77556 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636968456
transform 1 0 2300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636968456
transform 1 0 3404 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1
transform 1 0 4508 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1636968456
transform 1 0 4692 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1636968456
transform 1 0 5796 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636968456
transform 1 0 6900 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1636968456
transform 1 0 8004 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1
transform 1 0 9108 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1
transform 1 0 9660 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1636968456
transform 1 0 9844 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1636968456
transform 1 0 10948 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1636968456
transform 1 0 12052 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1636968456
transform 1 0 13156 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1
transform 1 0 14260 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1
transform 1 0 14812 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1636968456
transform 1 0 14996 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1636968456
transform 1 0 16100 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1636968456
transform 1 0 17204 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1636968456
transform 1 0 18308 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1
transform 1 0 19412 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1
transform 1 0 19964 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1636968456
transform 1 0 20148 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1636968456
transform 1 0 21252 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1636968456
transform 1 0 22356 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1636968456
transform 1 0 23460 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1
transform 1 0 24564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1
transform 1 0 25116 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1636968456
transform 1 0 25300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1636968456
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1636968456
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1636968456
transform 1 0 28612 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1
transform 1 0 29716 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1
transform 1 0 30268 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1636968456
transform 1 0 30452 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1636968456
transform 1 0 31556 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1636968456
transform 1 0 32660 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1636968456
transform 1 0 33764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1
transform 1 0 34868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1
transform 1 0 35420 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1636968456
transform 1 0 35604 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1636968456
transform 1 0 36708 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1636968456
transform 1 0 37812 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1636968456
transform 1 0 38916 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1
transform 1 0 40020 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1
transform 1 0 40572 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1636968456
transform 1 0 40756 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1636968456
transform 1 0 41860 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1636968456
transform 1 0 42964 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1636968456
transform 1 0 44068 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1
transform 1 0 45172 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1
transform 1 0 45724 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1636968456
transform 1 0 45908 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1636968456
transform 1 0 47012 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1636968456
transform 1 0 48116 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1636968456
transform 1 0 49220 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1
transform 1 0 50324 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1
transform 1 0 50876 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1636968456
transform 1 0 51060 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1636968456
transform 1 0 52164 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1636968456
transform 1 0 53268 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1636968456
transform 1 0 54372 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1
transform 1 0 55476 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1
transform 1 0 56028 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1636968456
transform 1 0 56212 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1636968456
transform 1 0 57316 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1636968456
transform 1 0 58420 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1636968456
transform 1 0 59524 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1
transform 1 0 60628 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1
transform 1 0 61180 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1636968456
transform 1 0 61364 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1636968456
transform 1 0 62468 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1636968456
transform 1 0 63572 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1636968456
transform 1 0 64676 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1
transform 1 0 65780 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1
transform 1 0 66332 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1636968456
transform 1 0 66516 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1636968456
transform 1 0 67620 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_725
timestamp 1636968456
transform 1 0 68724 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_737
timestamp 1636968456
transform 1 0 69828 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 1
transform 1 0 70932 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 1
transform 1 0 71484 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_757
timestamp 1636968456
transform 1 0 71668 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_769
timestamp 1636968456
transform 1 0 72772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_781
timestamp 1636968456
transform 1 0 73876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_793
timestamp 1636968456
transform 1 0 74980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 1
transform 1 0 76084 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 1
transform 1 0 76636 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_813
timestamp 1
transform 1 0 76820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_821
timestamp 1
transform 1 0 77556 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_6
timestamp 1636968456
transform 1 0 2576 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_18
timestamp 1636968456
transform 1 0 3680 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_30
timestamp 1636968456
transform 1 0 4784 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_42
timestamp 1636968456
transform 1 0 5888 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1
transform 1 0 6992 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636968456
transform 1 0 7268 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1636968456
transform 1 0 8372 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1636968456
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1636968456
transform 1 0 10580 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1
transform 1 0 11684 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1
transform 1 0 12236 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1636968456
transform 1 0 12420 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1636968456
transform 1 0 13524 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1636968456
transform 1 0 14628 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1636968456
transform 1 0 15732 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1
transform 1 0 16836 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1
transform 1 0 17388 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1636968456
transform 1 0 17572 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1636968456
transform 1 0 18676 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1636968456
transform 1 0 19780 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1636968456
transform 1 0 20884 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1
transform 1 0 21988 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1
transform 1 0 22540 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1636968456
transform 1 0 22724 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1636968456
transform 1 0 23828 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1636968456
transform 1 0 24932 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1636968456
transform 1 0 26036 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1
transform 1 0 27140 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1
transform 1 0 27692 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1636968456
transform 1 0 27876 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1636968456
transform 1 0 28980 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1636968456
transform 1 0 30084 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1636968456
transform 1 0 31188 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1
transform 1 0 32292 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1
transform 1 0 32844 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1636968456
transform 1 0 33028 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1636968456
transform 1 0 34132 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1636968456
transform 1 0 35236 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1636968456
transform 1 0 36340 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1
transform 1 0 37444 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1
transform 1 0 37996 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1636968456
transform 1 0 38180 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1636968456
transform 1 0 39284 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1636968456
transform 1 0 40388 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1636968456
transform 1 0 41492 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1
transform 1 0 42596 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1
transform 1 0 43148 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1636968456
transform 1 0 43332 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1636968456
transform 1 0 44436 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1636968456
transform 1 0 45540 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1636968456
transform 1 0 46644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1
transform 1 0 47748 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1
transform 1 0 48300 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1636968456
transform 1 0 48484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1636968456
transform 1 0 49588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1636968456
transform 1 0 50692 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1636968456
transform 1 0 51796 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1
transform 1 0 52900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1
transform 1 0 53452 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1636968456
transform 1 0 53636 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1636968456
transform 1 0 54740 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1636968456
transform 1 0 55844 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1636968456
transform 1 0 56948 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1
transform 1 0 58052 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1
transform 1 0 58604 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1636968456
transform 1 0 58788 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1636968456
transform 1 0 59892 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1636968456
transform 1 0 60996 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1636968456
transform 1 0 62100 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1
transform 1 0 63204 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1
transform 1 0 63756 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1636968456
transform 1 0 63940 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1636968456
transform 1 0 65044 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1636968456
transform 1 0 66148 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1636968456
transform 1 0 67252 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1
transform 1 0 68356 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1
transform 1 0 68908 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_729
timestamp 1636968456
transform 1 0 69092 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_741
timestamp 1636968456
transform 1 0 70196 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_753
timestamp 1636968456
transform 1 0 71300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_765
timestamp 1636968456
transform 1 0 72404 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 1
transform 1 0 73508 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 1
transform 1 0 74060 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_785
timestamp 1636968456
transform 1 0 74244 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_797
timestamp 1636968456
transform 1 0 75348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_809
timestamp 1636968456
transform 1 0 76452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_821
timestamp 1
transform 1 0 77556 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636968456
transform 1 0 2300 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1636968456
transform 1 0 3404 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1
transform 1 0 4508 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636968456
transform 1 0 4692 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1636968456
transform 1 0 5796 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1636968456
transform 1 0 6900 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1636968456
transform 1 0 8004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1
transform 1 0 9108 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1
transform 1 0 9660 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1636968456
transform 1 0 9844 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1636968456
transform 1 0 10948 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1636968456
transform 1 0 12052 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1636968456
transform 1 0 13156 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1
transform 1 0 14260 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1
transform 1 0 14812 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1636968456
transform 1 0 14996 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1636968456
transform 1 0 16100 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1636968456
transform 1 0 17204 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1636968456
transform 1 0 18308 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1
transform 1 0 19412 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1
transform 1 0 19964 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1636968456
transform 1 0 20148 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1636968456
transform 1 0 21252 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1636968456
transform 1 0 22356 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1636968456
transform 1 0 23460 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1
transform 1 0 24564 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1
transform 1 0 25116 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1636968456
transform 1 0 25300 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1636968456
transform 1 0 26404 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1636968456
transform 1 0 27508 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1636968456
transform 1 0 28612 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1
transform 1 0 29716 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1
transform 1 0 30268 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1636968456
transform 1 0 30452 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1636968456
transform 1 0 31556 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1636968456
transform 1 0 32660 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1636968456
transform 1 0 33764 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1
transform 1 0 34868 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1
transform 1 0 35420 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1636968456
transform 1 0 35604 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1636968456
transform 1 0 36708 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1636968456
transform 1 0 37812 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1636968456
transform 1 0 38916 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1
transform 1 0 40020 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1
transform 1 0 40572 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1636968456
transform 1 0 40756 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1636968456
transform 1 0 41860 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1636968456
transform 1 0 42964 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1636968456
transform 1 0 44068 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1
transform 1 0 45172 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1
transform 1 0 45724 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1636968456
transform 1 0 45908 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1636968456
transform 1 0 47012 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1636968456
transform 1 0 48116 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1636968456
transform 1 0 49220 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1
transform 1 0 50324 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1
transform 1 0 50876 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1636968456
transform 1 0 51060 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1636968456
transform 1 0 52164 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1636968456
transform 1 0 53268 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1636968456
transform 1 0 54372 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1
transform 1 0 55476 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1
transform 1 0 56028 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1636968456
transform 1 0 56212 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1636968456
transform 1 0 57316 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1636968456
transform 1 0 58420 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1636968456
transform 1 0 59524 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1
transform 1 0 60628 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1
transform 1 0 61180 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1636968456
transform 1 0 61364 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1636968456
transform 1 0 62468 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1636968456
transform 1 0 63572 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1636968456
transform 1 0 64676 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1
transform 1 0 65780 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1
transform 1 0 66332 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1636968456
transform 1 0 66516 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1636968456
transform 1 0 67620 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_725
timestamp 1636968456
transform 1 0 68724 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_737
timestamp 1636968456
transform 1 0 69828 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 1
transform 1 0 70932 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 1
transform 1 0 71484 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_757
timestamp 1636968456
transform 1 0 71668 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_769
timestamp 1636968456
transform 1 0 72772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_781
timestamp 1636968456
transform 1 0 73876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_793
timestamp 1636968456
transform 1 0 74980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 1
transform 1 0 76084 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 1
transform 1 0 76636 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_813
timestamp 1
transform 1 0 76820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_821
timestamp 1
transform 1 0 77556 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636968456
transform 1 0 2300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636968456
transform 1 0 3404 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1636968456
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636968456
transform 1 0 5612 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1
transform 1 0 6716 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1
transform 1 0 7084 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636968456
transform 1 0 7268 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1636968456
transform 1 0 8372 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1636968456
transform 1 0 9476 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1636968456
transform 1 0 10580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1
transform 1 0 11684 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1
transform 1 0 12236 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1636968456
transform 1 0 12420 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1636968456
transform 1 0 13524 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1636968456
transform 1 0 14628 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1636968456
transform 1 0 15732 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1
transform 1 0 16836 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1
transform 1 0 17388 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1636968456
transform 1 0 17572 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1636968456
transform 1 0 18676 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1636968456
transform 1 0 19780 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1636968456
transform 1 0 20884 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1
transform 1 0 21988 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1636968456
transform 1 0 22724 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1636968456
transform 1 0 23828 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1636968456
transform 1 0 24932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1636968456
transform 1 0 26036 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1
transform 1 0 27140 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1
transform 1 0 27692 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1636968456
transform 1 0 27876 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1636968456
transform 1 0 28980 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1636968456
transform 1 0 30084 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1636968456
transform 1 0 31188 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1
transform 1 0 32292 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1
transform 1 0 32844 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1636968456
transform 1 0 33028 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1636968456
transform 1 0 34132 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1636968456
transform 1 0 35236 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1636968456
transform 1 0 36340 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1
transform 1 0 37444 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1
transform 1 0 37996 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1636968456
transform 1 0 38180 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1636968456
transform 1 0 39284 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1636968456
transform 1 0 40388 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1636968456
transform 1 0 41492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1
transform 1 0 42596 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1
transform 1 0 43148 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1636968456
transform 1 0 43332 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1636968456
transform 1 0 44436 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1636968456
transform 1 0 45540 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1636968456
transform 1 0 46644 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1
transform 1 0 47748 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1
transform 1 0 48300 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1636968456
transform 1 0 48484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1636968456
transform 1 0 49588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1636968456
transform 1 0 50692 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1636968456
transform 1 0 51796 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1
transform 1 0 52900 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1
transform 1 0 53452 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1636968456
transform 1 0 53636 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1636968456
transform 1 0 54740 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1636968456
transform 1 0 55844 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1636968456
transform 1 0 56948 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1
transform 1 0 58052 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1
transform 1 0 58604 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1636968456
transform 1 0 58788 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1636968456
transform 1 0 59892 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1636968456
transform 1 0 60996 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1636968456
transform 1 0 62100 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1
transform 1 0 63204 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1
transform 1 0 63756 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1636968456
transform 1 0 63940 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1636968456
transform 1 0 65044 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1636968456
transform 1 0 66148 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1636968456
transform 1 0 67252 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1
transform 1 0 68356 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1
transform 1 0 68908 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_729
timestamp 1636968456
transform 1 0 69092 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_741
timestamp 1636968456
transform 1 0 70196 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_753
timestamp 1636968456
transform 1 0 71300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_765
timestamp 1636968456
transform 1 0 72404 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 1
transform 1 0 73508 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 1
transform 1 0 74060 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_785
timestamp 1636968456
transform 1 0 74244 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_797
timestamp 1636968456
transform 1 0 75348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_809
timestamp 1636968456
transform 1 0 76452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_821
timestamp 1
transform 1 0 77556 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636968456
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636968456
transform 1 0 3404 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1
transform 1 0 4508 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636968456
transform 1 0 4692 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636968456
transform 1 0 5796 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1636968456
transform 1 0 6900 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1636968456
transform 1 0 8004 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1
transform 1 0 9108 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1
transform 1 0 9660 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1636968456
transform 1 0 9844 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1636968456
transform 1 0 10948 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1636968456
transform 1 0 12052 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1636968456
transform 1 0 13156 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1
transform 1 0 14260 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1
transform 1 0 14812 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1636968456
transform 1 0 14996 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1636968456
transform 1 0 16100 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1636968456
transform 1 0 17204 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1636968456
transform 1 0 18308 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1
transform 1 0 19412 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1
transform 1 0 19964 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1636968456
transform 1 0 20148 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1636968456
transform 1 0 21252 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1636968456
transform 1 0 22356 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1636968456
transform 1 0 23460 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1
transform 1 0 24564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1
transform 1 0 25116 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1636968456
transform 1 0 25300 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1636968456
transform 1 0 26404 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1636968456
transform 1 0 27508 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1636968456
transform 1 0 28612 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1
transform 1 0 29716 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1
transform 1 0 30268 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1636968456
transform 1 0 30452 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1636968456
transform 1 0 31556 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1636968456
transform 1 0 32660 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1636968456
transform 1 0 33764 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1
transform 1 0 34868 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1
transform 1 0 35420 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1636968456
transform 1 0 35604 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1636968456
transform 1 0 36708 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1636968456
transform 1 0 37812 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1636968456
transform 1 0 38916 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1
transform 1 0 40020 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1
transform 1 0 40572 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1636968456
transform 1 0 40756 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1636968456
transform 1 0 41860 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1636968456
transform 1 0 42964 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1636968456
transform 1 0 44068 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1
transform 1 0 45172 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1
transform 1 0 45724 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1636968456
transform 1 0 45908 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1636968456
transform 1 0 47012 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1636968456
transform 1 0 48116 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1636968456
transform 1 0 49220 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1
transform 1 0 50324 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1
transform 1 0 50876 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1636968456
transform 1 0 51060 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1636968456
transform 1 0 52164 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1636968456
transform 1 0 53268 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1636968456
transform 1 0 54372 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1
transform 1 0 55476 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1
transform 1 0 56028 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1636968456
transform 1 0 56212 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1636968456
transform 1 0 57316 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1636968456
transform 1 0 58420 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1636968456
transform 1 0 59524 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1
transform 1 0 60628 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1
transform 1 0 61180 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1636968456
transform 1 0 61364 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1636968456
transform 1 0 62468 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1636968456
transform 1 0 63572 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1636968456
transform 1 0 64676 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1
transform 1 0 65780 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1
transform 1 0 66332 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1636968456
transform 1 0 66516 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1636968456
transform 1 0 67620 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_725
timestamp 1636968456
transform 1 0 68724 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_737
timestamp 1636968456
transform 1 0 69828 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 1
transform 1 0 70932 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 1
transform 1 0 71484 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_757
timestamp 1636968456
transform 1 0 71668 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_769
timestamp 1636968456
transform 1 0 72772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_781
timestamp 1636968456
transform 1 0 73876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_793
timestamp 1636968456
transform 1 0 74980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 1
transform 1 0 76084 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 1
transform 1 0 76636 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_813
timestamp 1
transform 1 0 76820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_821
timestamp 1
transform 1 0 77556 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636968456
transform 1 0 2300 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636968456
transform 1 0 3404 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1636968456
transform 1 0 4508 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1636968456
transform 1 0 5612 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1
transform 1 0 6716 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 7084 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636968456
transform 1 0 7268 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1636968456
transform 1 0 8372 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1636968456
transform 1 0 9476 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1636968456
transform 1 0 10580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1
transform 1 0 11684 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1
transform 1 0 12236 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1636968456
transform 1 0 12420 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1636968456
transform 1 0 13524 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1636968456
transform 1 0 14628 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1636968456
transform 1 0 15732 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1
transform 1 0 16836 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1
transform 1 0 17388 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1636968456
transform 1 0 17572 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1636968456
transform 1 0 18676 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1636968456
transform 1 0 19780 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1636968456
transform 1 0 20884 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1
transform 1 0 21988 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1
transform 1 0 22540 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636968456
transform 1 0 22724 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1636968456
transform 1 0 23828 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1636968456
transform 1 0 24932 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1636968456
transform 1 0 26036 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1
transform 1 0 27140 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1
transform 1 0 27692 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1636968456
transform 1 0 27876 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1636968456
transform 1 0 28980 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1636968456
transform 1 0 30084 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1636968456
transform 1 0 31188 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1
transform 1 0 32292 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1
transform 1 0 32844 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1636968456
transform 1 0 33028 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1636968456
transform 1 0 34132 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1636968456
transform 1 0 35236 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1636968456
transform 1 0 36340 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1
transform 1 0 37444 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1
transform 1 0 37996 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1636968456
transform 1 0 38180 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1636968456
transform 1 0 39284 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1636968456
transform 1 0 40388 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1636968456
transform 1 0 41492 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1
transform 1 0 42596 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1
transform 1 0 43148 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1636968456
transform 1 0 43332 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1636968456
transform 1 0 44436 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1636968456
transform 1 0 45540 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1636968456
transform 1 0 46644 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1
transform 1 0 47748 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1
transform 1 0 48300 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1636968456
transform 1 0 48484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1636968456
transform 1 0 49588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1636968456
transform 1 0 50692 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1636968456
transform 1 0 51796 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1
transform 1 0 52900 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1
transform 1 0 53452 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1636968456
transform 1 0 53636 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1636968456
transform 1 0 54740 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1636968456
transform 1 0 55844 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1636968456
transform 1 0 56948 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1
transform 1 0 58052 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1
transform 1 0 58604 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1636968456
transform 1 0 58788 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1636968456
transform 1 0 59892 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1636968456
transform 1 0 60996 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1636968456
transform 1 0 62100 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1
transform 1 0 63204 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1
transform 1 0 63756 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1636968456
transform 1 0 63940 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1636968456
transform 1 0 65044 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1636968456
transform 1 0 66148 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1636968456
transform 1 0 67252 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1
transform 1 0 68356 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1
transform 1 0 68908 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_729
timestamp 1636968456
transform 1 0 69092 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_741
timestamp 1636968456
transform 1 0 70196 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_753
timestamp 1636968456
transform 1 0 71300 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_765
timestamp 1636968456
transform 1 0 72404 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 1
transform 1 0 73508 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 1
transform 1 0 74060 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_785
timestamp 1636968456
transform 1 0 74244 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_797
timestamp 1636968456
transform 1 0 75348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_809
timestamp 1636968456
transform 1 0 76452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_821
timestamp 1
transform 1 0 77556 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_6
timestamp 1636968456
transform 1 0 2576 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_18
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1
transform 1 0 4416 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1636968456
transform 1 0 4692 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1636968456
transform 1 0 5796 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1636968456
transform 1 0 6900 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1636968456
transform 1 0 8004 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1
transform 1 0 9108 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1
transform 1 0 9660 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1636968456
transform 1 0 9844 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1636968456
transform 1 0 10948 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1636968456
transform 1 0 12052 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1636968456
transform 1 0 13156 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1
transform 1 0 14260 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1636968456
transform 1 0 14996 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1636968456
transform 1 0 16100 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1636968456
transform 1 0 17204 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1636968456
transform 1 0 18308 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1
transform 1 0 19412 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1
transform 1 0 19964 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1636968456
transform 1 0 20148 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1636968456
transform 1 0 21252 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1636968456
transform 1 0 22356 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1636968456
transform 1 0 23460 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1
transform 1 0 24564 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1
transform 1 0 25116 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1636968456
transform 1 0 25300 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1636968456
transform 1 0 26404 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1636968456
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1636968456
transform 1 0 28612 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1
transform 1 0 29716 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1
transform 1 0 30268 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1636968456
transform 1 0 30452 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1636968456
transform 1 0 31556 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1636968456
transform 1 0 32660 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1636968456
transform 1 0 33764 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1
transform 1 0 34868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1
transform 1 0 35420 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1636968456
transform 1 0 35604 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1636968456
transform 1 0 36708 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1636968456
transform 1 0 37812 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1636968456
transform 1 0 38916 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1
transform 1 0 40020 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1
transform 1 0 40572 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1636968456
transform 1 0 40756 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1636968456
transform 1 0 41860 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1636968456
transform 1 0 42964 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1636968456
transform 1 0 44068 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1
transform 1 0 45172 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1
transform 1 0 45724 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1636968456
transform 1 0 45908 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1636968456
transform 1 0 47012 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1636968456
transform 1 0 48116 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1636968456
transform 1 0 49220 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1
transform 1 0 50324 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1
transform 1 0 50876 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1636968456
transform 1 0 51060 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1636968456
transform 1 0 52164 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1636968456
transform 1 0 53268 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1636968456
transform 1 0 54372 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1
transform 1 0 55476 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1
transform 1 0 56028 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1636968456
transform 1 0 56212 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1636968456
transform 1 0 57316 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1636968456
transform 1 0 58420 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1636968456
transform 1 0 59524 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1
transform 1 0 60628 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1
transform 1 0 61180 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1636968456
transform 1 0 61364 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1636968456
transform 1 0 62468 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1636968456
transform 1 0 63572 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1636968456
transform 1 0 64676 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1
transform 1 0 65780 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1
transform 1 0 66332 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1636968456
transform 1 0 66516 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1636968456
transform 1 0 67620 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_725
timestamp 1636968456
transform 1 0 68724 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_737
timestamp 1636968456
transform 1 0 69828 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_749
timestamp 1
transform 1 0 70932 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_755
timestamp 1
transform 1 0 71484 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_757
timestamp 1636968456
transform 1 0 71668 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_769
timestamp 1636968456
transform 1 0 72772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_781
timestamp 1636968456
transform 1 0 73876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_793
timestamp 1636968456
transform 1 0 74980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_805
timestamp 1
transform 1 0 76084 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_811
timestamp 1
transform 1 0 76636 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_813
timestamp 1
transform 1 0 76820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_821
timestamp 1
transform 1 0 77556 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_6
timestamp 1636968456
transform 1 0 2576 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_18
timestamp 1636968456
transform 1 0 3680 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_30
timestamp 1636968456
transform 1 0 4784 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_42
timestamp 1636968456
transform 1 0 5888 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1
transform 1 0 6992 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1636968456
transform 1 0 7268 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1636968456
transform 1 0 8372 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1636968456
transform 1 0 9476 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1636968456
transform 1 0 10580 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1
transform 1 0 11684 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1
transform 1 0 12236 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1636968456
transform 1 0 12420 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1636968456
transform 1 0 13524 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1636968456
transform 1 0 14628 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1636968456
transform 1 0 15732 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1
transform 1 0 16836 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1
transform 1 0 17388 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636968456
transform 1 0 17572 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1636968456
transform 1 0 18676 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1636968456
transform 1 0 19780 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1636968456
transform 1 0 20884 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1
transform 1 0 21988 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1
transform 1 0 22540 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1636968456
transform 1 0 22724 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1636968456
transform 1 0 23828 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1636968456
transform 1 0 24932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1636968456
transform 1 0 26036 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1
transform 1 0 27140 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1
transform 1 0 27692 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1636968456
transform 1 0 27876 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1636968456
transform 1 0 28980 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1636968456
transform 1 0 30084 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1636968456
transform 1 0 31188 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1
transform 1 0 32292 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1
transform 1 0 32844 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1636968456
transform 1 0 33028 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1636968456
transform 1 0 34132 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1636968456
transform 1 0 35236 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1636968456
transform 1 0 36340 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1
transform 1 0 37444 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1
transform 1 0 37996 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1636968456
transform 1 0 38180 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1636968456
transform 1 0 39284 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1636968456
transform 1 0 40388 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1636968456
transform 1 0 41492 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1
transform 1 0 42596 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1
transform 1 0 43148 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1636968456
transform 1 0 43332 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1636968456
transform 1 0 44436 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1636968456
transform 1 0 45540 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1636968456
transform 1 0 46644 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1
transform 1 0 47748 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1
transform 1 0 48300 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1636968456
transform 1 0 48484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1636968456
transform 1 0 49588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1636968456
transform 1 0 50692 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1636968456
transform 1 0 51796 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1
transform 1 0 52900 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1
transform 1 0 53452 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1636968456
transform 1 0 53636 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1636968456
transform 1 0 54740 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1636968456
transform 1 0 55844 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1636968456
transform 1 0 56948 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1
transform 1 0 58052 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1
transform 1 0 58604 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1636968456
transform 1 0 58788 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1636968456
transform 1 0 59892 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1636968456
transform 1 0 60996 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1636968456
transform 1 0 62100 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1
transform 1 0 63204 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1
transform 1 0 63756 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1636968456
transform 1 0 63940 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1636968456
transform 1 0 65044 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1636968456
transform 1 0 66148 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1636968456
transform 1 0 67252 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1
transform 1 0 68356 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1
transform 1 0 68908 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_729
timestamp 1636968456
transform 1 0 69092 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_741
timestamp 1636968456
transform 1 0 70196 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_753
timestamp 1636968456
transform 1 0 71300 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_765
timestamp 1636968456
transform 1 0 72404 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_777
timestamp 1
transform 1 0 73508 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_783
timestamp 1
transform 1 0 74060 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_785
timestamp 1636968456
transform 1 0 74244 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_797
timestamp 1636968456
transform 1 0 75348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_809
timestamp 1636968456
transform 1 0 76452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_821
timestamp 1
transform 1 0 77556 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636968456
transform 1 0 2300 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636968456
transform 1 0 3404 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1
transform 1 0 4508 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636968456
transform 1 0 4692 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1636968456
transform 1 0 5796 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1636968456
transform 1 0 6900 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1636968456
transform 1 0 8004 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1
transform 1 0 9108 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1
transform 1 0 9660 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1636968456
transform 1 0 9844 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1636968456
transform 1 0 10948 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1636968456
transform 1 0 12052 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1636968456
transform 1 0 13156 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1
transform 1 0 14260 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1
transform 1 0 14812 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1636968456
transform 1 0 14996 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1636968456
transform 1 0 16100 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1636968456
transform 1 0 17204 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1636968456
transform 1 0 18308 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1
transform 1 0 19412 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1
transform 1 0 19964 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1636968456
transform 1 0 20148 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1636968456
transform 1 0 21252 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1636968456
transform 1 0 22356 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1636968456
transform 1 0 23460 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1
transform 1 0 24564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1
transform 1 0 25116 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1636968456
transform 1 0 25300 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1636968456
transform 1 0 26404 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1636968456
transform 1 0 27508 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1636968456
transform 1 0 28612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1
transform 1 0 29716 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1
transform 1 0 30268 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1636968456
transform 1 0 30452 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1636968456
transform 1 0 31556 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1636968456
transform 1 0 32660 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1636968456
transform 1 0 33764 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1
transform 1 0 34868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1
transform 1 0 35420 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1636968456
transform 1 0 35604 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1636968456
transform 1 0 36708 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1636968456
transform 1 0 37812 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1636968456
transform 1 0 38916 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1
transform 1 0 40020 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1
transform 1 0 40572 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1636968456
transform 1 0 40756 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1636968456
transform 1 0 41860 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1636968456
transform 1 0 42964 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1636968456
transform 1 0 44068 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1
transform 1 0 45172 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1
transform 1 0 45724 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1636968456
transform 1 0 45908 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1636968456
transform 1 0 47012 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1636968456
transform 1 0 48116 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1636968456
transform 1 0 49220 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1
transform 1 0 50324 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1
transform 1 0 50876 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1636968456
transform 1 0 51060 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1636968456
transform 1 0 52164 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1636968456
transform 1 0 53268 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1636968456
transform 1 0 54372 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1
transform 1 0 55476 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1
transform 1 0 56028 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1636968456
transform 1 0 56212 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1636968456
transform 1 0 57316 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1636968456
transform 1 0 58420 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1636968456
transform 1 0 59524 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1
transform 1 0 60628 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1
transform 1 0 61180 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1636968456
transform 1 0 61364 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1636968456
transform 1 0 62468 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1636968456
transform 1 0 63572 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1636968456
transform 1 0 64676 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1
transform 1 0 65780 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1
transform 1 0 66332 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1636968456
transform 1 0 66516 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1636968456
transform 1 0 67620 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_725
timestamp 1636968456
transform 1 0 68724 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_737
timestamp 1636968456
transform 1 0 69828 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_749
timestamp 1
transform 1 0 70932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_755
timestamp 1
transform 1 0 71484 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_757
timestamp 1636968456
transform 1 0 71668 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_769
timestamp 1636968456
transform 1 0 72772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_781
timestamp 1636968456
transform 1 0 73876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_793
timestamp 1636968456
transform 1 0 74980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_805
timestamp 1
transform 1 0 76084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_811
timestamp 1
transform 1 0 76636 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_813
timestamp 1
transform 1 0 76820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_821
timestamp 1
transform 1 0 77556 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_6
timestamp 1636968456
transform 1 0 2576 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_18
timestamp 1636968456
transform 1 0 3680 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_30
timestamp 1636968456
transform 1 0 4784 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_42
timestamp 1636968456
transform 1 0 5888 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp 1
transform 1 0 6992 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636968456
transform 1 0 7268 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1636968456
transform 1 0 8372 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1636968456
transform 1 0 9476 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1636968456
transform 1 0 10580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1
transform 1 0 11684 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1
transform 1 0 12236 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1636968456
transform 1 0 12420 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1636968456
transform 1 0 13524 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1636968456
transform 1 0 14628 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1636968456
transform 1 0 15732 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1
transform 1 0 16836 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1
transform 1 0 17388 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1636968456
transform 1 0 17572 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1636968456
transform 1 0 18676 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1636968456
transform 1 0 19780 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1636968456
transform 1 0 20884 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1
transform 1 0 21988 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1
transform 1 0 22540 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1636968456
transform 1 0 22724 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1636968456
transform 1 0 23828 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1636968456
transform 1 0 24932 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1636968456
transform 1 0 26036 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1
transform 1 0 27140 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1
transform 1 0 27692 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1636968456
transform 1 0 27876 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1636968456
transform 1 0 28980 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1636968456
transform 1 0 30084 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1636968456
transform 1 0 31188 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1
transform 1 0 32292 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1
transform 1 0 32844 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1636968456
transform 1 0 33028 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1636968456
transform 1 0 34132 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1636968456
transform 1 0 35236 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1636968456
transform 1 0 36340 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1
transform 1 0 37444 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1
transform 1 0 37996 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1636968456
transform 1 0 38180 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1636968456
transform 1 0 39284 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1636968456
transform 1 0 40388 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1636968456
transform 1 0 41492 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1
transform 1 0 42596 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1
transform 1 0 43148 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1636968456
transform 1 0 43332 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1636968456
transform 1 0 44436 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1636968456
transform 1 0 45540 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1636968456
transform 1 0 46644 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1
transform 1 0 47748 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1
transform 1 0 48300 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1636968456
transform 1 0 48484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1636968456
transform 1 0 49588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1636968456
transform 1 0 50692 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1636968456
transform 1 0 51796 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1
transform 1 0 52900 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1
transform 1 0 53452 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1636968456
transform 1 0 53636 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1636968456
transform 1 0 54740 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1636968456
transform 1 0 55844 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1636968456
transform 1 0 56948 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1
transform 1 0 58052 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1
transform 1 0 58604 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1636968456
transform 1 0 58788 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1636968456
transform 1 0 59892 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1636968456
transform 1 0 60996 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1636968456
transform 1 0 62100 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1
transform 1 0 63204 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1
transform 1 0 63756 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1636968456
transform 1 0 63940 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1636968456
transform 1 0 65044 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1636968456
transform 1 0 66148 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1636968456
transform 1 0 67252 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1
transform 1 0 68356 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1
transform 1 0 68908 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_729
timestamp 1636968456
transform 1 0 69092 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_741
timestamp 1636968456
transform 1 0 70196 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_753
timestamp 1636968456
transform 1 0 71300 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_765
timestamp 1636968456
transform 1 0 72404 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_777
timestamp 1
transform 1 0 73508 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_783
timestamp 1
transform 1 0 74060 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_785
timestamp 1636968456
transform 1 0 74244 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_797
timestamp 1636968456
transform 1 0 75348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_809
timestamp 1636968456
transform 1 0 76452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_821
timestamp 1
transform 1 0 77556 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636968456
transform 1 0 2300 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636968456
transform 1 0 3404 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 4508 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636968456
transform 1 0 4692 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636968456
transform 1 0 5796 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636968456
transform 1 0 6900 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1636968456
transform 1 0 8004 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1
transform 1 0 9108 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1
transform 1 0 9660 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1636968456
transform 1 0 9844 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1636968456
transform 1 0 10948 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1636968456
transform 1 0 12052 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1636968456
transform 1 0 13156 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1
transform 1 0 14260 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1
transform 1 0 14812 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1636968456
transform 1 0 14996 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1636968456
transform 1 0 16100 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1636968456
transform 1 0 17204 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1636968456
transform 1 0 18308 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1
transform 1 0 19412 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1
transform 1 0 19964 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1636968456
transform 1 0 20148 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1636968456
transform 1 0 21252 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1636968456
transform 1 0 22356 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1636968456
transform 1 0 23460 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1
transform 1 0 24564 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1
transform 1 0 25116 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1636968456
transform 1 0 25300 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1636968456
transform 1 0 26404 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1636968456
transform 1 0 27508 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1636968456
transform 1 0 28612 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1
transform 1 0 29716 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1
transform 1 0 30268 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1636968456
transform 1 0 30452 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1636968456
transform 1 0 31556 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1636968456
transform 1 0 32660 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1636968456
transform 1 0 33764 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1
transform 1 0 34868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1
transform 1 0 35420 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1636968456
transform 1 0 35604 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1636968456
transform 1 0 36708 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1636968456
transform 1 0 37812 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1636968456
transform 1 0 38916 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1
transform 1 0 40020 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1
transform 1 0 40572 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1636968456
transform 1 0 40756 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1636968456
transform 1 0 41860 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1636968456
transform 1 0 42964 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1636968456
transform 1 0 44068 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1
transform 1 0 45172 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1
transform 1 0 45724 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1636968456
transform 1 0 45908 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1636968456
transform 1 0 47012 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1636968456
transform 1 0 48116 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1636968456
transform 1 0 49220 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1
transform 1 0 50324 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1
transform 1 0 50876 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1636968456
transform 1 0 51060 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1636968456
transform 1 0 52164 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1636968456
transform 1 0 53268 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1636968456
transform 1 0 54372 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1
transform 1 0 55476 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1
transform 1 0 56028 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1636968456
transform 1 0 56212 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1636968456
transform 1 0 57316 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1636968456
transform 1 0 58420 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_625
timestamp 1636968456
transform 1 0 59524 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1
transform 1 0 60628 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1
transform 1 0 61180 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1636968456
transform 1 0 61364 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1636968456
transform 1 0 62468 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1636968456
transform 1 0 63572 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1636968456
transform 1 0 64676 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1
transform 1 0 65780 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1
transform 1 0 66332 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1636968456
transform 1 0 66516 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1636968456
transform 1 0 67620 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_725
timestamp 1636968456
transform 1 0 68724 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_737
timestamp 1636968456
transform 1 0 69828 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_749
timestamp 1
transform 1 0 70932 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_755
timestamp 1
transform 1 0 71484 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_757
timestamp 1636968456
transform 1 0 71668 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_769
timestamp 1636968456
transform 1 0 72772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_781
timestamp 1636968456
transform 1 0 73876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_793
timestamp 1636968456
transform 1 0 74980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_805
timestamp 1
transform 1 0 76084 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_811
timestamp 1
transform 1 0 76636 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_813
timestamp 1
transform 1 0 76820 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_821
timestamp 1
transform 1 0 77556 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_6
timestamp 1636968456
transform 1 0 2576 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_18
timestamp 1636968456
transform 1 0 3680 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_30
timestamp 1636968456
transform 1 0 4784 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_42
timestamp 1636968456
transform 1 0 5888 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1
transform 1 0 6992 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636968456
transform 1 0 7268 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1636968456
transform 1 0 8372 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1636968456
transform 1 0 9476 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1636968456
transform 1 0 10580 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1
transform 1 0 11684 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1
transform 1 0 12236 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1636968456
transform 1 0 12420 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1636968456
transform 1 0 13524 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1636968456
transform 1 0 14628 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1636968456
transform 1 0 15732 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1
transform 1 0 16836 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1
transform 1 0 17388 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1636968456
transform 1 0 17572 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1636968456
transform 1 0 18676 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1636968456
transform 1 0 19780 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1636968456
transform 1 0 20884 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1
transform 1 0 21988 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1636968456
transform 1 0 22724 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1636968456
transform 1 0 23828 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1636968456
transform 1 0 24932 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1636968456
transform 1 0 26036 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1
transform 1 0 27140 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1
transform 1 0 27692 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1636968456
transform 1 0 27876 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1636968456
transform 1 0 28980 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1636968456
transform 1 0 30084 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1636968456
transform 1 0 31188 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1
transform 1 0 32292 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1
transform 1 0 32844 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1636968456
transform 1 0 33028 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1636968456
transform 1 0 34132 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1636968456
transform 1 0 35236 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1636968456
transform 1 0 36340 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1
transform 1 0 37444 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1636968456
transform 1 0 38180 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1636968456
transform 1 0 39284 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1636968456
transform 1 0 40388 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1636968456
transform 1 0 41492 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1
transform 1 0 42596 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1
transform 1 0 43148 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1636968456
transform 1 0 43332 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1636968456
transform 1 0 44436 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1636968456
transform 1 0 45540 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1636968456
transform 1 0 46644 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1
transform 1 0 47748 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1
transform 1 0 48300 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1636968456
transform 1 0 48484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1636968456
transform 1 0 49588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1636968456
transform 1 0 50692 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1636968456
transform 1 0 51796 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1
transform 1 0 52900 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1
transform 1 0 53452 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1636968456
transform 1 0 53636 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1636968456
transform 1 0 54740 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1636968456
transform 1 0 55844 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1636968456
transform 1 0 56948 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1
transform 1 0 58052 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1
transform 1 0 58604 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1636968456
transform 1 0 58788 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1636968456
transform 1 0 59892 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1636968456
transform 1 0 60996 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1636968456
transform 1 0 62100 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1
transform 1 0 63204 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1
transform 1 0 63756 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1636968456
transform 1 0 63940 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1636968456
transform 1 0 65044 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1636968456
transform 1 0 66148 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1636968456
transform 1 0 67252 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1
transform 1 0 68356 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1
transform 1 0 68908 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_729
timestamp 1636968456
transform 1 0 69092 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_741
timestamp 1636968456
transform 1 0 70196 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_753
timestamp 1636968456
transform 1 0 71300 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_765
timestamp 1636968456
transform 1 0 72404 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_777
timestamp 1
transform 1 0 73508 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_783
timestamp 1
transform 1 0 74060 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_785
timestamp 1636968456
transform 1 0 74244 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_797
timestamp 1636968456
transform 1 0 75348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_809
timestamp 1636968456
transform 1 0 76452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_821
timestamp 1
transform 1 0 77556 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636968456
transform 1 0 2300 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1636968456
transform 1 0 3404 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1
transform 1 0 4508 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636968456
transform 1 0 4692 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1636968456
transform 1 0 5796 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1636968456
transform 1 0 6900 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1636968456
transform 1 0 8004 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1
transform 1 0 9108 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1
transform 1 0 9660 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1636968456
transform 1 0 9844 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1636968456
transform 1 0 10948 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1636968456
transform 1 0 12052 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1636968456
transform 1 0 13156 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1
transform 1 0 14260 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1
transform 1 0 14812 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1636968456
transform 1 0 14996 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1636968456
transform 1 0 16100 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1636968456
transform 1 0 17204 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1636968456
transform 1 0 18308 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1
transform 1 0 19412 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1
transform 1 0 19964 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1636968456
transform 1 0 20148 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1636968456
transform 1 0 21252 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1636968456
transform 1 0 22356 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1636968456
transform 1 0 23460 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1
transform 1 0 24564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1
transform 1 0 25116 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1636968456
transform 1 0 25300 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1636968456
transform 1 0 26404 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1636968456
transform 1 0 27508 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1636968456
transform 1 0 28612 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1
transform 1 0 29716 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1
transform 1 0 30268 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1636968456
transform 1 0 30452 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1636968456
transform 1 0 31556 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1636968456
transform 1 0 32660 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1636968456
transform 1 0 33764 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1
transform 1 0 34868 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1
transform 1 0 35420 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1636968456
transform 1 0 35604 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1636968456
transform 1 0 36708 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1636968456
transform 1 0 37812 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1636968456
transform 1 0 38916 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1
transform 1 0 40020 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1
transform 1 0 40572 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1636968456
transform 1 0 40756 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1636968456
transform 1 0 41860 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1636968456
transform 1 0 42964 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1636968456
transform 1 0 44068 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1
transform 1 0 45172 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1
transform 1 0 45724 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1636968456
transform 1 0 45908 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1636968456
transform 1 0 47012 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1636968456
transform 1 0 48116 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1636968456
transform 1 0 49220 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1
transform 1 0 50324 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1
transform 1 0 50876 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1636968456
transform 1 0 51060 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1636968456
transform 1 0 52164 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1636968456
transform 1 0 53268 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1636968456
transform 1 0 54372 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1
transform 1 0 55476 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1
transform 1 0 56028 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1636968456
transform 1 0 56212 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1636968456
transform 1 0 57316 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1636968456
transform 1 0 58420 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1636968456
transform 1 0 59524 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1
transform 1 0 60628 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1
transform 1 0 61180 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1636968456
transform 1 0 61364 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1636968456
transform 1 0 62468 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1636968456
transform 1 0 63572 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1636968456
transform 1 0 64676 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1
transform 1 0 65780 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1
transform 1 0 66332 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1636968456
transform 1 0 66516 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_713
timestamp 1636968456
transform 1 0 67620 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_725
timestamp 1636968456
transform 1 0 68724 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_737
timestamp 1636968456
transform 1 0 69828 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_749
timestamp 1
transform 1 0 70932 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_755
timestamp 1
transform 1 0 71484 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_757
timestamp 1636968456
transform 1 0 71668 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_769
timestamp 1636968456
transform 1 0 72772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_781
timestamp 1636968456
transform 1 0 73876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_793
timestamp 1636968456
transform 1 0 74980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_805
timestamp 1
transform 1 0 76084 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_811
timestamp 1
transform 1 0 76636 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_813
timestamp 1
transform 1 0 76820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_821
timestamp 1
transform 1 0 77556 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636968456
transform 1 0 2300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636968456
transform 1 0 3404 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1636968456
transform 1 0 4508 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1636968456
transform 1 0 5612 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1
transform 1 0 6716 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1
transform 1 0 7084 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1636968456
transform 1 0 7268 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1636968456
transform 1 0 8372 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1636968456
transform 1 0 9476 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1636968456
transform 1 0 10580 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1
transform 1 0 11684 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1
transform 1 0 12236 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1636968456
transform 1 0 12420 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1636968456
transform 1 0 13524 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1636968456
transform 1 0 14628 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1636968456
transform 1 0 15732 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1
transform 1 0 16836 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1636968456
transform 1 0 17572 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1636968456
transform 1 0 18676 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1636968456
transform 1 0 19780 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1636968456
transform 1 0 20884 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1
transform 1 0 21988 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1
transform 1 0 22540 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1636968456
transform 1 0 22724 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1636968456
transform 1 0 23828 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1636968456
transform 1 0 24932 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1636968456
transform 1 0 26036 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1
transform 1 0 27140 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1
transform 1 0 27692 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1636968456
transform 1 0 27876 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1636968456
transform 1 0 28980 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1636968456
transform 1 0 30084 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1636968456
transform 1 0 31188 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1
transform 1 0 32292 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1
transform 1 0 32844 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1636968456
transform 1 0 33028 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1636968456
transform 1 0 34132 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1636968456
transform 1 0 35236 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1636968456
transform 1 0 36340 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1
transform 1 0 37444 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1
transform 1 0 37996 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1636968456
transform 1 0 38180 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1636968456
transform 1 0 39284 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1636968456
transform 1 0 40388 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1636968456
transform 1 0 41492 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1
transform 1 0 42596 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1
transform 1 0 43148 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1636968456
transform 1 0 43332 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1636968456
transform 1 0 44436 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1636968456
transform 1 0 45540 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1636968456
transform 1 0 46644 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1
transform 1 0 47748 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1
transform 1 0 48300 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1636968456
transform 1 0 48484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1636968456
transform 1 0 49588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1636968456
transform 1 0 50692 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1636968456
transform 1 0 51796 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1
transform 1 0 52900 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1
transform 1 0 53452 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1636968456
transform 1 0 53636 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1636968456
transform 1 0 54740 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1636968456
transform 1 0 55844 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1636968456
transform 1 0 56948 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1
transform 1 0 58052 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1
transform 1 0 58604 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1636968456
transform 1 0 58788 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1636968456
transform 1 0 59892 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1636968456
transform 1 0 60996 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1636968456
transform 1 0 62100 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1
transform 1 0 63204 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1
transform 1 0 63756 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1636968456
transform 1 0 63940 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1636968456
transform 1 0 65044 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1636968456
transform 1 0 66148 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1636968456
transform 1 0 67252 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1
transform 1 0 68356 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1
transform 1 0 68908 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_729
timestamp 1636968456
transform 1 0 69092 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_741
timestamp 1636968456
transform 1 0 70196 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_753
timestamp 1636968456
transform 1 0 71300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_765
timestamp 1636968456
transform 1 0 72404 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_777
timestamp 1
transform 1 0 73508 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_783
timestamp 1
transform 1 0 74060 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_785
timestamp 1636968456
transform 1 0 74244 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_797
timestamp 1636968456
transform 1 0 75348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_809
timestamp 1636968456
transform 1 0 76452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_821
timestamp 1
transform 1 0 77556 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636968456
transform 1 0 2300 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636968456
transform 1 0 3404 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1
transform 1 0 4508 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636968456
transform 1 0 4692 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1636968456
transform 1 0 5796 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1636968456
transform 1 0 6900 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1636968456
transform 1 0 8004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1
transform 1 0 9108 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1
transform 1 0 9660 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1636968456
transform 1 0 9844 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1636968456
transform 1 0 10948 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1636968456
transform 1 0 12052 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1636968456
transform 1 0 13156 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1
transform 1 0 14260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1
transform 1 0 14812 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1636968456
transform 1 0 14996 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1636968456
transform 1 0 16100 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1636968456
transform 1 0 17204 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1636968456
transform 1 0 18308 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1
transform 1 0 19412 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1
transform 1 0 19964 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1636968456
transform 1 0 20148 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1636968456
transform 1 0 21252 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1636968456
transform 1 0 22356 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1636968456
transform 1 0 23460 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1
transform 1 0 24564 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1
transform 1 0 25116 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1636968456
transform 1 0 25300 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1636968456
transform 1 0 26404 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1636968456
transform 1 0 27508 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1636968456
transform 1 0 28612 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1
transform 1 0 29716 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1
transform 1 0 30268 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1636968456
transform 1 0 30452 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1636968456
transform 1 0 31556 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1636968456
transform 1 0 32660 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1636968456
transform 1 0 33764 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1
transform 1 0 34868 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1
transform 1 0 35420 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1636968456
transform 1 0 35604 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1636968456
transform 1 0 36708 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1636968456
transform 1 0 37812 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1636968456
transform 1 0 38916 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1
transform 1 0 40020 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1
transform 1 0 40572 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1636968456
transform 1 0 40756 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1636968456
transform 1 0 41860 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1636968456
transform 1 0 42964 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1636968456
transform 1 0 44068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1
transform 1 0 45172 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1
transform 1 0 45724 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1636968456
transform 1 0 45908 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1636968456
transform 1 0 47012 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1636968456
transform 1 0 48116 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1636968456
transform 1 0 49220 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1
transform 1 0 50324 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1
transform 1 0 50876 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1636968456
transform 1 0 51060 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1636968456
transform 1 0 52164 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1636968456
transform 1 0 53268 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1636968456
transform 1 0 54372 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1
transform 1 0 55476 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1
transform 1 0 56028 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1636968456
transform 1 0 56212 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1636968456
transform 1 0 57316 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1636968456
transform 1 0 58420 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_625
timestamp 1636968456
transform 1 0 59524 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1
transform 1 0 60628 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1
transform 1 0 61180 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1636968456
transform 1 0 61364 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1636968456
transform 1 0 62468 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1636968456
transform 1 0 63572 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1636968456
transform 1 0 64676 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1
transform 1 0 65780 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1
transform 1 0 66332 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1636968456
transform 1 0 66516 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1636968456
transform 1 0 67620 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_725
timestamp 1636968456
transform 1 0 68724 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_737
timestamp 1636968456
transform 1 0 69828 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_749
timestamp 1
transform 1 0 70932 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_755
timestamp 1
transform 1 0 71484 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_757
timestamp 1636968456
transform 1 0 71668 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_769
timestamp 1636968456
transform 1 0 72772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_781
timestamp 1636968456
transform 1 0 73876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_793
timestamp 1636968456
transform 1 0 74980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_805
timestamp 1
transform 1 0 76084 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_811
timestamp 1
transform 1 0 76636 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_813
timestamp 1
transform 1 0 76820 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_821
timestamp 1
transform 1 0 77556 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636968456
transform 1 0 2300 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636968456
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636968456
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1636968456
transform 1 0 5612 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1
transform 1 0 6716 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1
transform 1 0 7084 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1636968456
transform 1 0 7268 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1636968456
transform 1 0 8372 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1636968456
transform 1 0 9476 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1636968456
transform 1 0 10580 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1
transform 1 0 11684 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1
transform 1 0 12236 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1636968456
transform 1 0 12420 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1636968456
transform 1 0 13524 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1636968456
transform 1 0 14628 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1636968456
transform 1 0 15732 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1
transform 1 0 16836 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1
transform 1 0 17388 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1636968456
transform 1 0 17572 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1636968456
transform 1 0 18676 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1636968456
transform 1 0 19780 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1636968456
transform 1 0 20884 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1
transform 1 0 21988 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1
transform 1 0 22540 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1636968456
transform 1 0 22724 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1636968456
transform 1 0 23828 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1636968456
transform 1 0 24932 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1636968456
transform 1 0 26036 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1
transform 1 0 27140 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1
transform 1 0 27692 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1636968456
transform 1 0 27876 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1636968456
transform 1 0 28980 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1636968456
transform 1 0 30084 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1636968456
transform 1 0 31188 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1
transform 1 0 32292 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1
transform 1 0 32844 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1636968456
transform 1 0 33028 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1636968456
transform 1 0 34132 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1636968456
transform 1 0 35236 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1636968456
transform 1 0 36340 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1
transform 1 0 37444 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1
transform 1 0 37996 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1636968456
transform 1 0 38180 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1636968456
transform 1 0 39284 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1636968456
transform 1 0 40388 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1636968456
transform 1 0 41492 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1
transform 1 0 42596 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1
transform 1 0 43148 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1636968456
transform 1 0 43332 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1636968456
transform 1 0 44436 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1636968456
transform 1 0 45540 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1636968456
transform 1 0 46644 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1
transform 1 0 47748 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1
transform 1 0 48300 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1636968456
transform 1 0 48484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1636968456
transform 1 0 49588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1636968456
transform 1 0 50692 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1636968456
transform 1 0 51796 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1
transform 1 0 52900 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1
transform 1 0 53452 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1636968456
transform 1 0 53636 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1636968456
transform 1 0 54740 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1636968456
transform 1 0 55844 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1636968456
transform 1 0 56948 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1
transform 1 0 58052 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1
transform 1 0 58604 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1636968456
transform 1 0 58788 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_629
timestamp 1636968456
transform 1 0 59892 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_641
timestamp 1636968456
transform 1 0 60996 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_653
timestamp 1636968456
transform 1 0 62100 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1
transform 1 0 63204 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1
transform 1 0 63756 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1636968456
transform 1 0 63940 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1636968456
transform 1 0 65044 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1636968456
transform 1 0 66148 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1636968456
transform 1 0 67252 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1
transform 1 0 68356 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1
transform 1 0 68908 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_729
timestamp 1636968456
transform 1 0 69092 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_741
timestamp 1636968456
transform 1 0 70196 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_753
timestamp 1636968456
transform 1 0 71300 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_765
timestamp 1636968456
transform 1 0 72404 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_777
timestamp 1
transform 1 0 73508 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_783
timestamp 1
transform 1 0 74060 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_785
timestamp 1636968456
transform 1 0 74244 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_797
timestamp 1636968456
transform 1 0 75348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_809
timestamp 1636968456
transform 1 0 76452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_821
timestamp 1
transform 1 0 77556 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636968456
transform 1 0 2300 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636968456
transform 1 0 3404 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1
transform 1 0 4508 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1636968456
transform 1 0 4692 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1636968456
transform 1 0 5796 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1636968456
transform 1 0 6900 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1636968456
transform 1 0 8004 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1
transform 1 0 9108 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1
transform 1 0 9660 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1636968456
transform 1 0 9844 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1636968456
transform 1 0 10948 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1636968456
transform 1 0 12052 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1636968456
transform 1 0 13156 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1
transform 1 0 14260 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1
transform 1 0 14812 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1636968456
transform 1 0 14996 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1636968456
transform 1 0 16100 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1636968456
transform 1 0 17204 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1636968456
transform 1 0 18308 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1
transform 1 0 19412 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1
transform 1 0 19964 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1636968456
transform 1 0 20148 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1636968456
transform 1 0 21252 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1636968456
transform 1 0 22356 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1636968456
transform 1 0 23460 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1
transform 1 0 24564 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1
transform 1 0 25116 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1636968456
transform 1 0 25300 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1636968456
transform 1 0 26404 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1636968456
transform 1 0 27508 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1636968456
transform 1 0 28612 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1
transform 1 0 29716 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1
transform 1 0 30268 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1636968456
transform 1 0 30452 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1636968456
transform 1 0 31556 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1636968456
transform 1 0 32660 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1636968456
transform 1 0 33764 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1
transform 1 0 34868 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1
transform 1 0 35420 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1636968456
transform 1 0 35604 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1636968456
transform 1 0 36708 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1636968456
transform 1 0 37812 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1636968456
transform 1 0 38916 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1
transform 1 0 40020 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1
transform 1 0 40572 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1636968456
transform 1 0 40756 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1636968456
transform 1 0 41860 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1636968456
transform 1 0 42964 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1636968456
transform 1 0 44068 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1
transform 1 0 45172 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1
transform 1 0 45724 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1636968456
transform 1 0 45908 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1636968456
transform 1 0 47012 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1636968456
transform 1 0 48116 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1636968456
transform 1 0 49220 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1
transform 1 0 50324 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1
transform 1 0 50876 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1636968456
transform 1 0 51060 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1636968456
transform 1 0 52164 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1636968456
transform 1 0 53268 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1636968456
transform 1 0 54372 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1
transform 1 0 55476 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1
transform 1 0 56028 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1636968456
transform 1 0 56212 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1636968456
transform 1 0 57316 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1636968456
transform 1 0 58420 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_625
timestamp 1636968456
transform 1 0 59524 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1
transform 1 0 60628 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1
transform 1 0 61180 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1636968456
transform 1 0 61364 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1636968456
transform 1 0 62468 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1636968456
transform 1 0 63572 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1636968456
transform 1 0 64676 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1
transform 1 0 65780 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1
transform 1 0 66332 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_701
timestamp 1636968456
transform 1 0 66516 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_713
timestamp 1636968456
transform 1 0 67620 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_725
timestamp 1636968456
transform 1 0 68724 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_737
timestamp 1636968456
transform 1 0 69828 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_749
timestamp 1
transform 1 0 70932 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_755
timestamp 1
transform 1 0 71484 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_757
timestamp 1636968456
transform 1 0 71668 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_769
timestamp 1636968456
transform 1 0 72772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_781
timestamp 1636968456
transform 1 0 73876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_793
timestamp 1636968456
transform 1 0 74980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_805
timestamp 1
transform 1 0 76084 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_811
timestamp 1
transform 1 0 76636 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_813
timestamp 1
transform 1 0 76820 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_821
timestamp 1
transform 1 0 77556 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_6
timestamp 1636968456
transform 1 0 2576 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_18
timestamp 1636968456
transform 1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_30
timestamp 1636968456
transform 1 0 4784 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_42
timestamp 1636968456
transform 1 0 5888 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 1
transform 1 0 6992 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1636968456
transform 1 0 7268 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1636968456
transform 1 0 8372 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1636968456
transform 1 0 9476 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1636968456
transform 1 0 10580 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1
transform 1 0 11684 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1
transform 1 0 12236 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1636968456
transform 1 0 12420 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1636968456
transform 1 0 13524 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1636968456
transform 1 0 14628 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1636968456
transform 1 0 15732 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1
transform 1 0 16836 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1
transform 1 0 17388 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1636968456
transform 1 0 17572 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1636968456
transform 1 0 18676 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1636968456
transform 1 0 19780 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1636968456
transform 1 0 20884 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1
transform 1 0 21988 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1
transform 1 0 22540 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1636968456
transform 1 0 22724 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1636968456
transform 1 0 23828 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1636968456
transform 1 0 24932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1636968456
transform 1 0 26036 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1
transform 1 0 27140 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1
transform 1 0 27692 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1636968456
transform 1 0 27876 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1636968456
transform 1 0 28980 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1636968456
transform 1 0 30084 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1636968456
transform 1 0 31188 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1
transform 1 0 32292 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1
transform 1 0 32844 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1636968456
transform 1 0 33028 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1636968456
transform 1 0 34132 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1636968456
transform 1 0 35236 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1636968456
transform 1 0 36340 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1
transform 1 0 37444 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1
transform 1 0 37996 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1636968456
transform 1 0 38180 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1636968456
transform 1 0 39284 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1636968456
transform 1 0 40388 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1636968456
transform 1 0 41492 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1
transform 1 0 42596 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1
transform 1 0 43148 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1636968456
transform 1 0 43332 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1636968456
transform 1 0 44436 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1636968456
transform 1 0 45540 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1636968456
transform 1 0 46644 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1
transform 1 0 47748 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1
transform 1 0 48300 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1636968456
transform 1 0 48484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1636968456
transform 1 0 49588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1636968456
transform 1 0 50692 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1636968456
transform 1 0 51796 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1
transform 1 0 52900 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1
transform 1 0 53452 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1636968456
transform 1 0 53636 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1636968456
transform 1 0 54740 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1636968456
transform 1 0 55844 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1636968456
transform 1 0 56948 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1
transform 1 0 58052 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1
transform 1 0 58604 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1636968456
transform 1 0 58788 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1636968456
transform 1 0 59892 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1636968456
transform 1 0 60996 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_653
timestamp 1636968456
transform 1 0 62100 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1
transform 1 0 63204 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1
transform 1 0 63756 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1636968456
transform 1 0 63940 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1636968456
transform 1 0 65044 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_697
timestamp 1636968456
transform 1 0 66148 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_709
timestamp 1636968456
transform 1 0 67252 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 1
transform 1 0 68356 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 1
transform 1 0 68908 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_729
timestamp 1636968456
transform 1 0 69092 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_741
timestamp 1636968456
transform 1 0 70196 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_753
timestamp 1636968456
transform 1 0 71300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_765
timestamp 1636968456
transform 1 0 72404 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_777
timestamp 1
transform 1 0 73508 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_783
timestamp 1
transform 1 0 74060 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_785
timestamp 1636968456
transform 1 0 74244 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_797
timestamp 1636968456
transform 1 0 75348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_809
timestamp 1636968456
transform 1 0 76452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_821
timestamp 1
transform 1 0 77556 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636968456
transform 1 0 2300 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636968456
transform 1 0 3404 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1
transform 1 0 4508 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636968456
transform 1 0 4692 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1636968456
transform 1 0 5796 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1636968456
transform 1 0 6900 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1636968456
transform 1 0 8004 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1
transform 1 0 9108 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1
transform 1 0 9660 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1636968456
transform 1 0 9844 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1636968456
transform 1 0 10948 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1636968456
transform 1 0 12052 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1636968456
transform 1 0 13156 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1
transform 1 0 14260 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1
transform 1 0 14812 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1636968456
transform 1 0 14996 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1636968456
transform 1 0 16100 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1636968456
transform 1 0 17204 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1636968456
transform 1 0 18308 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1
transform 1 0 19412 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1
transform 1 0 19964 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1636968456
transform 1 0 20148 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1636968456
transform 1 0 21252 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1636968456
transform 1 0 22356 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1636968456
transform 1 0 23460 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1
transform 1 0 24564 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1
transform 1 0 25116 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1636968456
transform 1 0 25300 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1636968456
transform 1 0 26404 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1636968456
transform 1 0 27508 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1636968456
transform 1 0 28612 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1
transform 1 0 29716 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1
transform 1 0 30268 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1636968456
transform 1 0 30452 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1636968456
transform 1 0 31556 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1636968456
transform 1 0 32660 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1636968456
transform 1 0 33764 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1
transform 1 0 34868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1
transform 1 0 35420 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1636968456
transform 1 0 35604 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1636968456
transform 1 0 36708 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1636968456
transform 1 0 37812 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1636968456
transform 1 0 38916 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1
transform 1 0 40020 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1
transform 1 0 40572 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1636968456
transform 1 0 40756 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1636968456
transform 1 0 41860 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1636968456
transform 1 0 42964 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1636968456
transform 1 0 44068 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1
transform 1 0 45172 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1
transform 1 0 45724 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1636968456
transform 1 0 45908 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1636968456
transform 1 0 47012 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1636968456
transform 1 0 48116 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1636968456
transform 1 0 49220 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1
transform 1 0 50324 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1
transform 1 0 50876 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1636968456
transform 1 0 51060 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1636968456
transform 1 0 52164 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1636968456
transform 1 0 53268 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1636968456
transform 1 0 54372 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1
transform 1 0 55476 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1
transform 1 0 56028 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1636968456
transform 1 0 56212 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1636968456
transform 1 0 57316 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1636968456
transform 1 0 58420 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1636968456
transform 1 0 59524 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1
transform 1 0 60628 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1
transform 1 0 61180 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1636968456
transform 1 0 61364 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_657
timestamp 1636968456
transform 1 0 62468 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_669
timestamp 1636968456
transform 1 0 63572 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_681
timestamp 1636968456
transform 1 0 64676 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1
transform 1 0 65780 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1
transform 1 0 66332 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1636968456
transform 1 0 66516 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_713
timestamp 1636968456
transform 1 0 67620 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_725
timestamp 1636968456
transform 1 0 68724 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_737
timestamp 1636968456
transform 1 0 69828 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_749
timestamp 1
transform 1 0 70932 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_755
timestamp 1
transform 1 0 71484 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_757
timestamp 1636968456
transform 1 0 71668 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_769
timestamp 1636968456
transform 1 0 72772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_781
timestamp 1636968456
transform 1 0 73876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_793
timestamp 1636968456
transform 1 0 74980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_805
timestamp 1
transform 1 0 76084 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_811
timestamp 1
transform 1 0 76636 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_813
timestamp 1
transform 1 0 76820 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_821
timestamp 1
transform 1 0 77556 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636968456
transform 1 0 2300 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636968456
transform 1 0 3404 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1636968456
transform 1 0 4508 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1636968456
transform 1 0 5612 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1
transform 1 0 6716 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1
transform 1 0 7084 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1636968456
transform 1 0 7268 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1636968456
transform 1 0 8372 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1636968456
transform 1 0 9476 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1636968456
transform 1 0 10580 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1
transform 1 0 11684 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1
transform 1 0 12236 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1636968456
transform 1 0 12420 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1636968456
transform 1 0 13524 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1636968456
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1636968456
transform 1 0 15732 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1
transform 1 0 16836 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1
transform 1 0 17388 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1636968456
transform 1 0 17572 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1636968456
transform 1 0 18676 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1636968456
transform 1 0 19780 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1636968456
transform 1 0 20884 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1
transform 1 0 21988 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1
transform 1 0 22540 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1636968456
transform 1 0 22724 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1636968456
transform 1 0 23828 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1636968456
transform 1 0 24932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1636968456
transform 1 0 26036 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1
transform 1 0 27140 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1
transform 1 0 27692 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1636968456
transform 1 0 27876 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1636968456
transform 1 0 28980 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1636968456
transform 1 0 30084 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1636968456
transform 1 0 31188 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1
transform 1 0 32292 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1
transform 1 0 32844 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1636968456
transform 1 0 33028 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1636968456
transform 1 0 34132 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1636968456
transform 1 0 35236 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1636968456
transform 1 0 36340 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1
transform 1 0 37444 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1
transform 1 0 37996 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1636968456
transform 1 0 38180 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1636968456
transform 1 0 39284 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1636968456
transform 1 0 40388 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1636968456
transform 1 0 41492 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1
transform 1 0 42596 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1
transform 1 0 43148 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1636968456
transform 1 0 43332 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1636968456
transform 1 0 44436 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1636968456
transform 1 0 45540 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1636968456
transform 1 0 46644 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1
transform 1 0 47748 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1
transform 1 0 48300 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1636968456
transform 1 0 48484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1636968456
transform 1 0 49588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1636968456
transform 1 0 50692 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1636968456
transform 1 0 51796 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1
transform 1 0 52900 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1
transform 1 0 53452 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1636968456
transform 1 0 53636 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1636968456
transform 1 0 54740 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1636968456
transform 1 0 55844 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1636968456
transform 1 0 56948 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1
transform 1 0 58052 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1
transform 1 0 58604 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1636968456
transform 1 0 58788 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1636968456
transform 1 0 59892 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1636968456
transform 1 0 60996 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_653
timestamp 1636968456
transform 1 0 62100 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1
transform 1 0 63204 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1
transform 1 0 63756 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1636968456
transform 1 0 63940 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1636968456
transform 1 0 65044 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_697
timestamp 1
transform 1 0 66148 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_703
timestamp 1
transform 1 0 66700 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_707
timestamp 1636968456
transform 1 0 67068 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_719
timestamp 1
transform 1 0 68172 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1
transform 1 0 68908 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_729
timestamp 1636968456
transform 1 0 69092 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_741
timestamp 1636968456
transform 1 0 70196 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_753
timestamp 1636968456
transform 1 0 71300 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_765
timestamp 1636968456
transform 1 0 72404 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_777
timestamp 1
transform 1 0 73508 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_783
timestamp 1
transform 1 0 74060 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_785
timestamp 1636968456
transform 1 0 74244 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_797
timestamp 1636968456
transform 1 0 75348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_809
timestamp 1636968456
transform 1 0 76452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_821
timestamp 1
transform 1 0 77556 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636968456
transform 1 0 2300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636968456
transform 1 0 3404 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1
transform 1 0 4508 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636968456
transform 1 0 4692 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1636968456
transform 1 0 5796 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1636968456
transform 1 0 6900 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1636968456
transform 1 0 8004 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1
transform 1 0 9108 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1
transform 1 0 9660 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1636968456
transform 1 0 9844 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1636968456
transform 1 0 10948 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1636968456
transform 1 0 12052 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1636968456
transform 1 0 13156 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1
transform 1 0 14260 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1
transform 1 0 14812 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1636968456
transform 1 0 14996 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1636968456
transform 1 0 16100 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1636968456
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1636968456
transform 1 0 18308 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1
transform 1 0 19412 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1
transform 1 0 19964 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1636968456
transform 1 0 20148 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1636968456
transform 1 0 21252 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1636968456
transform 1 0 22356 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1636968456
transform 1 0 23460 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1
transform 1 0 24564 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1
transform 1 0 25116 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1636968456
transform 1 0 25300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1636968456
transform 1 0 26404 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1636968456
transform 1 0 27508 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1636968456
transform 1 0 28612 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1
transform 1 0 29716 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1
transform 1 0 30268 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1636968456
transform 1 0 30452 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1636968456
transform 1 0 31556 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1636968456
transform 1 0 32660 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1636968456
transform 1 0 33764 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1
transform 1 0 34868 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1
transform 1 0 35420 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1636968456
transform 1 0 35604 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1636968456
transform 1 0 36708 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1636968456
transform 1 0 37812 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1636968456
transform 1 0 38916 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1
transform 1 0 40020 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1
transform 1 0 40572 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1636968456
transform 1 0 40756 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1636968456
transform 1 0 41860 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1636968456
transform 1 0 42964 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1636968456
transform 1 0 44068 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1
transform 1 0 45172 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1
transform 1 0 45724 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1636968456
transform 1 0 45908 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1636968456
transform 1 0 47012 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1636968456
transform 1 0 48116 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1636968456
transform 1 0 49220 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1
transform 1 0 50324 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1
transform 1 0 50876 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1636968456
transform 1 0 51060 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1636968456
transform 1 0 52164 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1636968456
transform 1 0 53268 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1636968456
transform 1 0 54372 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1
transform 1 0 55476 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1
transform 1 0 56028 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1636968456
transform 1 0 56212 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1636968456
transform 1 0 57316 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1636968456
transform 1 0 58420 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1636968456
transform 1 0 59524 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1
transform 1 0 60628 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1
transform 1 0 61180 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1636968456
transform 1 0 61364 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1636968456
transform 1 0 62468 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1636968456
transform 1 0 63572 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1636968456
transform 1 0 64676 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1
transform 1 0 65780 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1
transform 1 0 66332 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_721
timestamp 1636968456
transform 1 0 68356 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_733
timestamp 1636968456
transform 1 0 69460 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_745
timestamp 1
transform 1 0 70564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_751
timestamp 1
transform 1 0 71116 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_755
timestamp 1
transform 1 0 71484 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_757
timestamp 1636968456
transform 1 0 71668 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_769
timestamp 1636968456
transform 1 0 72772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_781
timestamp 1636968456
transform 1 0 73876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_793
timestamp 1636968456
transform 1 0 74980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_805
timestamp 1
transform 1 0 76084 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_811
timestamp 1
transform 1 0 76636 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_813
timestamp 1
transform 1 0 76820 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_821
timestamp 1
transform 1 0 77556 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636968456
transform 1 0 2300 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636968456
transform 1 0 3404 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636968456
transform 1 0 4508 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1636968456
transform 1 0 5612 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1
transform 1 0 6716 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1
transform 1 0 7084 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1636968456
transform 1 0 7268 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1636968456
transform 1 0 8372 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1636968456
transform 1 0 9476 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1636968456
transform 1 0 10580 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1
transform 1 0 11684 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1
transform 1 0 12236 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1636968456
transform 1 0 12420 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1636968456
transform 1 0 13524 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1636968456
transform 1 0 14628 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1636968456
transform 1 0 15732 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1
transform 1 0 16836 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1
transform 1 0 17388 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1636968456
transform 1 0 17572 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1636968456
transform 1 0 18676 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1636968456
transform 1 0 19780 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1636968456
transform 1 0 20884 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1
transform 1 0 21988 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1
transform 1 0 22540 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1636968456
transform 1 0 22724 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1636968456
transform 1 0 23828 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1636968456
transform 1 0 24932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1636968456
transform 1 0 26036 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1
transform 1 0 27140 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1
transform 1 0 27692 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1636968456
transform 1 0 27876 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1636968456
transform 1 0 28980 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1636968456
transform 1 0 30084 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1636968456
transform 1 0 31188 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1
transform 1 0 32292 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1636968456
transform 1 0 33028 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1636968456
transform 1 0 34132 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1636968456
transform 1 0 35236 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1636968456
transform 1 0 36340 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1
transform 1 0 37444 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1
transform 1 0 37996 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1636968456
transform 1 0 38180 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1636968456
transform 1 0 39284 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1636968456
transform 1 0 40388 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1636968456
transform 1 0 41492 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1
transform 1 0 42596 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1
transform 1 0 43148 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1636968456
transform 1 0 43332 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1636968456
transform 1 0 44436 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1636968456
transform 1 0 45540 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1636968456
transform 1 0 46644 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1
transform 1 0 47748 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1
transform 1 0 48300 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1636968456
transform 1 0 48484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1636968456
transform 1 0 49588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1636968456
transform 1 0 50692 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1636968456
transform 1 0 51796 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1
transform 1 0 52900 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1
transform 1 0 53452 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1636968456
transform 1 0 53636 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1636968456
transform 1 0 54740 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1636968456
transform 1 0 55844 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1636968456
transform 1 0 56948 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1
transform 1 0 58052 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1
transform 1 0 58604 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1636968456
transform 1 0 58788 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1636968456
transform 1 0 59892 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1636968456
transform 1 0 60996 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1636968456
transform 1 0 62100 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1
transform 1 0 63204 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1
transform 1 0 63756 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1636968456
transform 1 0 63940 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_685
timestamp 1
transform 1 0 65044 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_691
timestamp 1
transform 1 0 65596 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_707
timestamp 1636968456
transform 1 0 67068 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_719
timestamp 1
transform 1 0 68172 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1
transform 1 0 68908 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_729
timestamp 1
transform 1 0 69092 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_763
timestamp 1636968456
transform 1 0 72220 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_775
timestamp 1
transform 1 0 73324 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_783
timestamp 1
transform 1 0 74060 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_785
timestamp 1636968456
transform 1 0 74244 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_797
timestamp 1636968456
transform 1 0 75348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_809
timestamp 1
transform 1 0 76452 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_817
timestamp 1
transform 1 0 77188 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636968456
transform 1 0 2300 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1636968456
transform 1 0 3404 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1
transform 1 0 4508 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636968456
transform 1 0 4692 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1636968456
transform 1 0 5796 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1636968456
transform 1 0 6900 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1636968456
transform 1 0 8004 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1
transform 1 0 9108 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1
transform 1 0 9660 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1636968456
transform 1 0 9844 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1636968456
transform 1 0 10948 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1636968456
transform 1 0 12052 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1636968456
transform 1 0 13156 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1
transform 1 0 14260 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1
transform 1 0 14812 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1636968456
transform 1 0 14996 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1636968456
transform 1 0 16100 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1636968456
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1636968456
transform 1 0 18308 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1
transform 1 0 19412 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1
transform 1 0 19964 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1636968456
transform 1 0 20148 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1636968456
transform 1 0 21252 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1636968456
transform 1 0 22356 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1636968456
transform 1 0 23460 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1
transform 1 0 24564 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1
transform 1 0 25116 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1636968456
transform 1 0 25300 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1636968456
transform 1 0 26404 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1636968456
transform 1 0 27508 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1636968456
transform 1 0 28612 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1
transform 1 0 29716 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1
transform 1 0 30268 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1636968456
transform 1 0 30452 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1636968456
transform 1 0 31556 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1636968456
transform 1 0 32660 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1636968456
transform 1 0 33764 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1
transform 1 0 34868 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1
transform 1 0 35420 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1636968456
transform 1 0 35604 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1636968456
transform 1 0 36708 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1636968456
transform 1 0 37812 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1636968456
transform 1 0 38916 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1
transform 1 0 40020 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1
transform 1 0 40572 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1636968456
transform 1 0 40756 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1636968456
transform 1 0 41860 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1636968456
transform 1 0 42964 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1636968456
transform 1 0 44068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1
transform 1 0 45172 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1
transform 1 0 45724 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1636968456
transform 1 0 45908 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1636968456
transform 1 0 47012 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1636968456
transform 1 0 48116 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1636968456
transform 1 0 49220 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1
transform 1 0 50324 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1
transform 1 0 50876 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1636968456
transform 1 0 51060 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1636968456
transform 1 0 52164 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1636968456
transform 1 0 53268 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1636968456
transform 1 0 54372 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1
transform 1 0 55476 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1
transform 1 0 56028 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_589
timestamp 1
transform 1 0 56212 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1636968456
transform 1 0 58420 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_625
timestamp 1636968456
transform 1 0 59524 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1
transform 1 0 60628 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1
transform 1 0 61180 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_645
timestamp 1636968456
transform 1 0 61364 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_657
timestamp 1636968456
transform 1 0 62468 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_669
timestamp 1636968456
transform 1 0 63572 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_681
timestamp 1636968456
transform 1 0 64676 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1
transform 1 0 65780 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1
transform 1 0 66332 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_701
timestamp 1636968456
transform 1 0 66516 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_713
timestamp 1636968456
transform 1 0 67620 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_725
timestamp 1636968456
transform 1 0 68724 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_737
timestamp 1
transform 1 0 69828 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_750
timestamp 1
transform 1 0 71024 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_757
timestamp 1636968456
transform 1 0 71668 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_769
timestamp 1636968456
transform 1 0 72772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_781
timestamp 1636968456
transform 1 0 73876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_793
timestamp 1636968456
transform 1 0 74980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_805
timestamp 1
transform 1 0 76084 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_811
timestamp 1
transform 1 0 76636 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_813
timestamp 1
transform 1 0 76820 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_821
timestamp 1
transform 1 0 77556 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_6
timestamp 1636968456
transform 1 0 2576 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_18
timestamp 1636968456
transform 1 0 3680 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_30
timestamp 1636968456
transform 1 0 4784 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_42
timestamp 1636968456
transform 1 0 5888 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1
transform 1 0 6992 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636968456
transform 1 0 7268 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1636968456
transform 1 0 8372 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1636968456
transform 1 0 9476 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1636968456
transform 1 0 10580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1
transform 1 0 11684 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1
transform 1 0 12236 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1636968456
transform 1 0 12420 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1636968456
transform 1 0 13524 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1636968456
transform 1 0 14628 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1636968456
transform 1 0 15732 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1
transform 1 0 16836 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1
transform 1 0 17388 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1636968456
transform 1 0 17572 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1636968456
transform 1 0 18676 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1636968456
transform 1 0 19780 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1636968456
transform 1 0 20884 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1
transform 1 0 21988 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1
transform 1 0 22540 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1636968456
transform 1 0 22724 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1636968456
transform 1 0 23828 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1636968456
transform 1 0 24932 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1636968456
transform 1 0 26036 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1
transform 1 0 27140 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1
transform 1 0 27692 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1636968456
transform 1 0 27876 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1636968456
transform 1 0 28980 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1636968456
transform 1 0 30084 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1636968456
transform 1 0 31188 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1
transform 1 0 32292 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1
transform 1 0 32844 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1636968456
transform 1 0 33028 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1636968456
transform 1 0 34132 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1636968456
transform 1 0 35236 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1636968456
transform 1 0 36340 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1
transform 1 0 37444 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1
transform 1 0 37996 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1636968456
transform 1 0 38180 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1636968456
transform 1 0 39284 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1636968456
transform 1 0 40388 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1636968456
transform 1 0 41492 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1
transform 1 0 42596 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1
transform 1 0 43148 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1636968456
transform 1 0 43332 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1636968456
transform 1 0 44436 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1636968456
transform 1 0 45540 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1636968456
transform 1 0 46644 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1
transform 1 0 47748 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1
transform 1 0 48300 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1636968456
transform 1 0 48484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1636968456
transform 1 0 49588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1636968456
transform 1 0 50692 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1636968456
transform 1 0 51796 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1
transform 1 0 52900 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1
transform 1 0 53452 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1636968456
transform 1 0 53636 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1636968456
transform 1 0 54740 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_585
timestamp 1
transform 1 0 55844 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_589
timestamp 1
transform 1 0 56212 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_597
timestamp 1
transform 1 0 56948 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_601
timestamp 1
transform 1 0 57316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_610
timestamp 1
transform 1 0 58144 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_617
timestamp 1636968456
transform 1 0 58788 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_629
timestamp 1
transform 1 0 59892 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_633
timestamp 1
transform 1 0 60260 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_657
timestamp 1636968456
transform 1 0 62468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_669
timestamp 1
transform 1 0 63572 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_673
timestamp 1636968456
transform 1 0 63940 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_685
timestamp 1636968456
transform 1 0 65044 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_697
timestamp 1636968456
transform 1 0 66148 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_709
timestamp 1636968456
transform 1 0 67252 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1
transform 1 0 68356 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1
transform 1 0 68908 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_729
timestamp 1
transform 1 0 69092 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_737
timestamp 1
transform 1 0 69828 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_760
timestamp 1636968456
transform 1 0 71944 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_772
timestamp 1636968456
transform 1 0 73048 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_785
timestamp 1
transform 1 0 74244 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_794
timestamp 1636968456
transform 1 0 75072 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_806
timestamp 1636968456
transform 1 0 76176 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_818
timestamp 1
transform 1 0 77280 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636968456
transform 1 0 2300 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636968456
transform 1 0 3404 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1
transform 1 0 4508 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636968456
transform 1 0 4692 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1636968456
transform 1 0 5796 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1636968456
transform 1 0 6900 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1636968456
transform 1 0 8004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1
transform 1 0 9108 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1
transform 1 0 9660 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1636968456
transform 1 0 9844 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1636968456
transform 1 0 10948 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1636968456
transform 1 0 12052 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1636968456
transform 1 0 13156 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1
transform 1 0 14260 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1
transform 1 0 14812 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1636968456
transform 1 0 14996 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1636968456
transform 1 0 16100 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1636968456
transform 1 0 17204 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1636968456
transform 1 0 18308 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1
transform 1 0 19412 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1
transform 1 0 19964 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1636968456
transform 1 0 20148 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1636968456
transform 1 0 21252 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1636968456
transform 1 0 22356 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1636968456
transform 1 0 23460 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1
transform 1 0 24564 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1
transform 1 0 25116 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1636968456
transform 1 0 25300 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1636968456
transform 1 0 26404 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1636968456
transform 1 0 27508 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1636968456
transform 1 0 28612 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1
transform 1 0 29716 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1
transform 1 0 30268 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1636968456
transform 1 0 30452 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1636968456
transform 1 0 31556 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1636968456
transform 1 0 32660 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1636968456
transform 1 0 33764 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1
transform 1 0 34868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1
transform 1 0 35420 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1636968456
transform 1 0 35604 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1636968456
transform 1 0 36708 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1636968456
transform 1 0 37812 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1636968456
transform 1 0 38916 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1
transform 1 0 40020 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1
transform 1 0 40572 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1636968456
transform 1 0 40756 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1636968456
transform 1 0 41860 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1636968456
transform 1 0 42964 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1636968456
transform 1 0 44068 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1
transform 1 0 45172 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1
transform 1 0 45724 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1636968456
transform 1 0 45908 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1636968456
transform 1 0 47012 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1636968456
transform 1 0 48116 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1636968456
transform 1 0 49220 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1
transform 1 0 50324 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1
transform 1 0 50876 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1636968456
transform 1 0 51060 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1636968456
transform 1 0 52164 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1636968456
transform 1 0 53268 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1636968456
transform 1 0 54372 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1
transform 1 0 55476 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1
transform 1 0 56028 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1636968456
transform 1 0 56212 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1636968456
transform 1 0 57316 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1636968456
transform 1 0 58420 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_625
timestamp 1
transform 1 0 59524 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_642
timestamp 1
transform 1 0 61088 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_645
timestamp 1636968456
transform 1 0 61364 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_657
timestamp 1636968456
transform 1 0 62468 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_669
timestamp 1636968456
transform 1 0 63572 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_681
timestamp 1636968456
transform 1 0 64676 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1
transform 1 0 65780 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1
transform 1 0 66332 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_704
timestamp 1636968456
transform 1 0 66792 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_716
timestamp 1636968456
transform 1 0 67896 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_728
timestamp 1636968456
transform 1 0 69000 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_740
timestamp 1
transform 1 0 70104 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_744
timestamp 1
transform 1 0 70472 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_749
timestamp 1
transform 1 0 70932 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_755
timestamp 1
transform 1 0 71484 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_757
timestamp 1
transform 1 0 71668 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_765
timestamp 1
transform 1 0 72404 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_774
timestamp 1
transform 1 0 73232 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_782
timestamp 1
transform 1 0 73968 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_810
timestamp 1
transform 1 0 76544 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_813
timestamp 1
transform 1 0 76820 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_821
timestamp 1
transform 1 0 77556 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636968456
transform 1 0 2300 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636968456
transform 1 0 3404 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1636968456
transform 1 0 4508 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1636968456
transform 1 0 5612 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1
transform 1 0 6716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1636968456
transform 1 0 7268 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1636968456
transform 1 0 8372 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1636968456
transform 1 0 9476 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1636968456
transform 1 0 10580 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1
transform 1 0 11684 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1
transform 1 0 12236 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1636968456
transform 1 0 12420 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1636968456
transform 1 0 13524 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1636968456
transform 1 0 14628 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1636968456
transform 1 0 15732 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1
transform 1 0 16836 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1
transform 1 0 17388 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1636968456
transform 1 0 17572 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1636968456
transform 1 0 18676 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1636968456
transform 1 0 19780 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1636968456
transform 1 0 20884 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1
transform 1 0 21988 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1
transform 1 0 22540 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1636968456
transform 1 0 22724 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1636968456
transform 1 0 23828 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1636968456
transform 1 0 24932 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1636968456
transform 1 0 26036 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1
transform 1 0 27140 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1
transform 1 0 27692 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1636968456
transform 1 0 27876 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1636968456
transform 1 0 28980 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1636968456
transform 1 0 30084 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1636968456
transform 1 0 31188 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1
transform 1 0 32292 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1
transform 1 0 32844 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1636968456
transform 1 0 33028 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1636968456
transform 1 0 34132 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1636968456
transform 1 0 35236 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1636968456
transform 1 0 36340 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1
transform 1 0 37444 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1
transform 1 0 37996 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1636968456
transform 1 0 38180 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1636968456
transform 1 0 39284 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1636968456
transform 1 0 40388 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1636968456
transform 1 0 41492 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1
transform 1 0 42596 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1
transform 1 0 43148 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1636968456
transform 1 0 43332 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1636968456
transform 1 0 44436 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1636968456
transform 1 0 45540 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1636968456
transform 1 0 46644 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1
transform 1 0 47748 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1
transform 1 0 48300 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1636968456
transform 1 0 48484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1636968456
transform 1 0 49588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1636968456
transform 1 0 50692 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1636968456
transform 1 0 51796 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1
transform 1 0 52900 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1
transform 1 0 53452 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1636968456
transform 1 0 53636 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1636968456
transform 1 0 54740 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1636968456
transform 1 0 55844 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1636968456
transform 1 0 56948 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1
transform 1 0 58052 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1
transform 1 0 58604 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_617
timestamp 1636968456
transform 1 0 58788 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_629
timestamp 1
transform 1 0 59892 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_639
timestamp 1636968456
transform 1 0 60812 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_651
timestamp 1636968456
transform 1 0 61916 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_663
timestamp 1
transform 1 0 63020 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1
transform 1 0 63756 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_673
timestamp 1636968456
transform 1 0 63940 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_685
timestamp 1
transform 1 0 65044 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_698
timestamp 1636968456
transform 1 0 66240 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_710
timestamp 1636968456
transform 1 0 67344 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_722
timestamp 1
transform 1 0 68448 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_729
timestamp 1636968456
transform 1 0 69092 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_741
timestamp 1636968456
transform 1 0 70196 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_753
timestamp 1636968456
transform 1 0 71300 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_765
timestamp 1636968456
transform 1 0 72404 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_777
timestamp 1
transform 1 0 73508 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_783
timestamp 1
transform 1 0 74060 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_785
timestamp 1636968456
transform 1 0 74244 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_797
timestamp 1636968456
transform 1 0 75348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_809
timestamp 1636968456
transform 1 0 76452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_821
timestamp 1
transform 1 0 77556 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1636968456
transform 1 0 2300 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1636968456
transform 1 0 3404 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1
transform 1 0 4508 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636968456
transform 1 0 4692 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1636968456
transform 1 0 5796 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1636968456
transform 1 0 6900 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1636968456
transform 1 0 8004 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1
transform 1 0 9108 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1
transform 1 0 9660 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1636968456
transform 1 0 9844 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1636968456
transform 1 0 10948 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1636968456
transform 1 0 12052 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1636968456
transform 1 0 13156 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1
transform 1 0 14260 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1
transform 1 0 14812 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1636968456
transform 1 0 14996 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1636968456
transform 1 0 16100 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1636968456
transform 1 0 17204 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1636968456
transform 1 0 18308 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1
transform 1 0 19412 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1636968456
transform 1 0 20148 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1636968456
transform 1 0 21252 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1636968456
transform 1 0 22356 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1636968456
transform 1 0 23460 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1
transform 1 0 24564 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1
transform 1 0 25116 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1636968456
transform 1 0 25300 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1636968456
transform 1 0 26404 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1636968456
transform 1 0 27508 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1636968456
transform 1 0 28612 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1
transform 1 0 29716 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1
transform 1 0 30268 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1636968456
transform 1 0 30452 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1636968456
transform 1 0 31556 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1636968456
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1636968456
transform 1 0 33764 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1
transform 1 0 34868 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1
transform 1 0 35420 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1636968456
transform 1 0 35604 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1636968456
transform 1 0 36708 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1636968456
transform 1 0 37812 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1636968456
transform 1 0 38916 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1
transform 1 0 40020 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1
transform 1 0 40572 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1636968456
transform 1 0 40756 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1636968456
transform 1 0 41860 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1636968456
transform 1 0 42964 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1636968456
transform 1 0 44068 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1
transform 1 0 45172 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1
transform 1 0 45724 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1636968456
transform 1 0 45908 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1636968456
transform 1 0 47012 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1636968456
transform 1 0 48116 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1636968456
transform 1 0 49220 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1
transform 1 0 50324 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1
transform 1 0 50876 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1636968456
transform 1 0 51060 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1636968456
transform 1 0 52164 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1636968456
transform 1 0 53268 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1636968456
transform 1 0 54372 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1
transform 1 0 55476 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1
transform 1 0 56028 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1636968456
transform 1 0 56212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_601
timestamp 1
transform 1 0 57316 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_606
timestamp 1636968456
transform 1 0 57776 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_618
timestamp 1636968456
transform 1 0 58880 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_630
timestamp 1636968456
transform 1 0 59984 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_642
timestamp 1
transform 1 0 61088 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_645
timestamp 1636968456
transform 1 0 61364 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_657
timestamp 1636968456
transform 1 0 62468 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_669
timestamp 1
transform 1 0 63572 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_697
timestamp 1
transform 1 0 66148 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_709
timestamp 1636968456
transform 1 0 67252 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_721
timestamp 1636968456
transform 1 0 68356 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_733
timestamp 1636968456
transform 1 0 69460 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_745
timestamp 1
transform 1 0 70564 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_753
timestamp 1
transform 1 0 71300 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_757
timestamp 1636968456
transform 1 0 71668 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_769
timestamp 1636968456
transform 1 0 72772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_781
timestamp 1636968456
transform 1 0 73876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_793
timestamp 1
transform 1 0 74980 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_798
timestamp 1636968456
transform 1 0 75440 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_810
timestamp 1
transform 1 0 76544 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_813
timestamp 1
transform 1 0 76820 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_817
timestamp 1
transform 1 0 77188 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1636968456
transform 1 0 2300 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1636968456
transform 1 0 3404 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1636968456
transform 1 0 4508 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1636968456
transform 1 0 5612 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1
transform 1 0 6716 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1
transform 1 0 7084 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1636968456
transform 1 0 7268 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1636968456
transform 1 0 8372 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1636968456
transform 1 0 9476 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1636968456
transform 1 0 10580 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1
transform 1 0 11684 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1
transform 1 0 12236 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1636968456
transform 1 0 12420 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1636968456
transform 1 0 13524 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1636968456
transform 1 0 14628 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1636968456
transform 1 0 15732 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1
transform 1 0 16836 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1
transform 1 0 17388 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1636968456
transform 1 0 17572 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1636968456
transform 1 0 18676 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1636968456
transform 1 0 19780 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1636968456
transform 1 0 20884 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1
transform 1 0 21988 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1
transform 1 0 22540 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1636968456
transform 1 0 22724 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1636968456
transform 1 0 23828 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1636968456
transform 1 0 24932 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1636968456
transform 1 0 26036 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1
transform 1 0 27140 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1
transform 1 0 27692 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1636968456
transform 1 0 27876 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1636968456
transform 1 0 28980 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1636968456
transform 1 0 30084 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1636968456
transform 1 0 31188 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1
transform 1 0 32292 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1
transform 1 0 32844 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1636968456
transform 1 0 33028 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1636968456
transform 1 0 34132 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1636968456
transform 1 0 35236 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1636968456
transform 1 0 36340 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1
transform 1 0 37444 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1
transform 1 0 37996 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1636968456
transform 1 0 38180 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1636968456
transform 1 0 39284 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1636968456
transform 1 0 40388 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1636968456
transform 1 0 41492 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1
transform 1 0 42596 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1
transform 1 0 43148 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1636968456
transform 1 0 43332 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1636968456
transform 1 0 44436 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1636968456
transform 1 0 45540 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1636968456
transform 1 0 46644 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1
transform 1 0 47748 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1
transform 1 0 48300 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1636968456
transform 1 0 48484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1636968456
transform 1 0 49588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1636968456
transform 1 0 50692 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1636968456
transform 1 0 51796 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1
transform 1 0 52900 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1
transform 1 0 53452 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1636968456
transform 1 0 53636 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1636968456
transform 1 0 54740 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1636968456
transform 1 0 55844 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1636968456
transform 1 0 56948 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1
transform 1 0 58052 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1
transform 1 0 58604 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_617
timestamp 1636968456
transform 1 0 58788 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_629
timestamp 1636968456
transform 1 0 59892 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_641
timestamp 1636968456
transform 1 0 60996 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_653
timestamp 1636968456
transform 1 0 62100 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1
transform 1 0 63204 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_671
timestamp 1
transform 1 0 63756 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_673
timestamp 1636968456
transform 1 0 63940 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_685
timestamp 1636968456
transform 1 0 65044 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_697
timestamp 1636968456
transform 1 0 66148 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_709
timestamp 1
transform 1 0 67252 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_721
timestamp 1
transform 1 0 68356 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_727
timestamp 1
transform 1 0 68908 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_729
timestamp 1636968456
transform 1 0 69092 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_741
timestamp 1636968456
transform 1 0 70196 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_753
timestamp 1636968456
transform 1 0 71300 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_765
timestamp 1636968456
transform 1 0 72404 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_777
timestamp 1
transform 1 0 73508 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_783
timestamp 1
transform 1 0 74060 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_785
timestamp 1636968456
transform 1 0 74244 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_797
timestamp 1636968456
transform 1 0 75348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_809
timestamp 1
transform 1 0 76452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_817
timestamp 1
transform 1 0 77188 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1636968456
transform 1 0 2300 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1636968456
transform 1 0 3404 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1
transform 1 0 4508 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1636968456
transform 1 0 4692 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1636968456
transform 1 0 5796 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1636968456
transform 1 0 6900 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1636968456
transform 1 0 8004 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1
transform 1 0 9108 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1
transform 1 0 9660 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1636968456
transform 1 0 9844 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1636968456
transform 1 0 10948 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1636968456
transform 1 0 12052 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1636968456
transform 1 0 13156 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1
transform 1 0 14260 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1
transform 1 0 14812 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1636968456
transform 1 0 14996 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1636968456
transform 1 0 16100 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1636968456
transform 1 0 17204 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1636968456
transform 1 0 18308 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1
transform 1 0 19412 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1
transform 1 0 19964 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1636968456
transform 1 0 20148 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1636968456
transform 1 0 21252 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1636968456
transform 1 0 22356 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1636968456
transform 1 0 23460 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1
transform 1 0 24564 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1
transform 1 0 25116 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1636968456
transform 1 0 25300 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1636968456
transform 1 0 26404 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1636968456
transform 1 0 27508 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1636968456
transform 1 0 28612 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1
transform 1 0 29716 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1
transform 1 0 30268 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1636968456
transform 1 0 30452 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1636968456
transform 1 0 31556 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1636968456
transform 1 0 32660 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1636968456
transform 1 0 33764 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1
transform 1 0 34868 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1
transform 1 0 35420 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1636968456
transform 1 0 35604 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1636968456
transform 1 0 36708 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1636968456
transform 1 0 37812 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1636968456
transform 1 0 38916 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1
transform 1 0 40020 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1
transform 1 0 40572 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1636968456
transform 1 0 40756 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1636968456
transform 1 0 41860 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1636968456
transform 1 0 42964 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1636968456
transform 1 0 44068 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1
transform 1 0 45172 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1
transform 1 0 45724 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1636968456
transform 1 0 45908 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1636968456
transform 1 0 47012 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1636968456
transform 1 0 48116 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1636968456
transform 1 0 49220 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1
transform 1 0 50324 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1
transform 1 0 50876 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1636968456
transform 1 0 51060 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1636968456
transform 1 0 52164 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1636968456
transform 1 0 53268 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1636968456
transform 1 0 54372 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1
transform 1 0 55476 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1
transform 1 0 56028 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_589
timestamp 1
transform 1 0 56212 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_597
timestamp 1
transform 1 0 56948 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_603
timestamp 1
transform 1 0 57500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_609
timestamp 1636968456
transform 1 0 58052 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_621
timestamp 1636968456
transform 1 0 59156 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_633
timestamp 1
transform 1 0 60260 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_641
timestamp 1
transform 1 0 60996 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_645
timestamp 1636968456
transform 1 0 61364 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_657
timestamp 1
transform 1 0 62468 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_661
timestamp 1
transform 1 0 62836 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_682
timestamp 1636968456
transform 1 0 64768 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_694
timestamp 1
transform 1 0 65872 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_701
timestamp 1636968456
transform 1 0 66516 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_713
timestamp 1
transform 1 0 67620 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_735
timestamp 1636968456
transform 1 0 69644 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_747
timestamp 1
transform 1 0 70748 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_755
timestamp 1
transform 1 0 71484 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_757
timestamp 1636968456
transform 1 0 71668 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_769
timestamp 1636968456
transform 1 0 72772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_781
timestamp 1
transform 1 0 73876 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_792
timestamp 1636968456
transform 1 0 74888 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_804
timestamp 1
transform 1 0 75992 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_808
timestamp 1
transform 1 0 76360 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_813
timestamp 1
transform 1 0 76820 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_817
timestamp 1
transform 1 0 77188 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1636968456
transform 1 0 2300 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1636968456
transform 1 0 3404 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1636968456
transform 1 0 4508 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1636968456
transform 1 0 5612 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1
transform 1 0 6716 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1
transform 1 0 7084 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1636968456
transform 1 0 7268 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1636968456
transform 1 0 8372 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1636968456
transform 1 0 9476 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1636968456
transform 1 0 10580 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1
transform 1 0 11684 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1
transform 1 0 12236 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1636968456
transform 1 0 12420 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1636968456
transform 1 0 13524 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1636968456
transform 1 0 14628 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1636968456
transform 1 0 15732 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1
transform 1 0 16836 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1
transform 1 0 17388 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1636968456
transform 1 0 17572 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1636968456
transform 1 0 18676 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1636968456
transform 1 0 19780 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1636968456
transform 1 0 20884 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1
transform 1 0 21988 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1
transform 1 0 22540 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1636968456
transform 1 0 22724 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1636968456
transform 1 0 23828 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1636968456
transform 1 0 24932 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1636968456
transform 1 0 26036 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1
transform 1 0 27140 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1
transform 1 0 27692 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1636968456
transform 1 0 27876 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1636968456
transform 1 0 28980 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1636968456
transform 1 0 30084 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1636968456
transform 1 0 31188 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1
transform 1 0 32292 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1
transform 1 0 32844 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1636968456
transform 1 0 33028 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1636968456
transform 1 0 34132 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1636968456
transform 1 0 35236 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1636968456
transform 1 0 36340 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1
transform 1 0 37444 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1
transform 1 0 37996 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1636968456
transform 1 0 38180 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1636968456
transform 1 0 39284 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1636968456
transform 1 0 40388 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1636968456
transform 1 0 41492 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1
transform 1 0 42596 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1
transform 1 0 43148 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1636968456
transform 1 0 43332 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1636968456
transform 1 0 44436 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1636968456
transform 1 0 45540 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1636968456
transform 1 0 46644 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1
transform 1 0 47748 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1
transform 1 0 48300 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1636968456
transform 1 0 48484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1636968456
transform 1 0 49588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1636968456
transform 1 0 50692 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1636968456
transform 1 0 51796 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1
transform 1 0 52900 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1
transform 1 0 53452 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1636968456
transform 1 0 53636 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1636968456
transform 1 0 54740 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1636968456
transform 1 0 55844 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1636968456
transform 1 0 56948 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1
transform 1 0 58052 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1
transform 1 0 58604 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_617
timestamp 1636968456
transform 1 0 58788 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_629
timestamp 1636968456
transform 1 0 59892 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_641
timestamp 1636968456
transform 1 0 60996 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_653
timestamp 1636968456
transform 1 0 62100 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1
transform 1 0 63204 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1
transform 1 0 63756 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_673
timestamp 1636968456
transform 1 0 63940 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_685
timestamp 1
transform 1 0 65044 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_709
timestamp 1636968456
transform 1 0 67252 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_721
timestamp 1
transform 1 0 68356 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_727
timestamp 1
transform 1 0 68908 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_729
timestamp 1636968456
transform 1 0 69092 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_741
timestamp 1
transform 1 0 70196 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_747
timestamp 1
transform 1 0 70748 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_761
timestamp 1636968456
transform 1 0 72036 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_773
timestamp 1
transform 1 0 73140 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_781
timestamp 1
transform 1 0 73876 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_785
timestamp 1
transform 1 0 74244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_793
timestamp 1
transform 1 0 74980 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_804
timestamp 1636968456
transform 1 0 75992 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_816
timestamp 1
transform 1 0 77096 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636968456
transform 1 0 2300 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636968456
transform 1 0 3404 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1
transform 1 0 4508 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636968456
transform 1 0 4692 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1636968456
transform 1 0 5796 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1636968456
transform 1 0 6900 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1636968456
transform 1 0 8004 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1
transform 1 0 9108 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1
transform 1 0 9660 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1636968456
transform 1 0 9844 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1636968456
transform 1 0 10948 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1636968456
transform 1 0 12052 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1636968456
transform 1 0 13156 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1
transform 1 0 14260 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1
transform 1 0 14812 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1636968456
transform 1 0 14996 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1636968456
transform 1 0 16100 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1636968456
transform 1 0 17204 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1636968456
transform 1 0 18308 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1
transform 1 0 19412 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1
transform 1 0 19964 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1636968456
transform 1 0 20148 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1636968456
transform 1 0 21252 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1636968456
transform 1 0 22356 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1636968456
transform 1 0 23460 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1
transform 1 0 24564 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1
transform 1 0 25116 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1636968456
transform 1 0 25300 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1636968456
transform 1 0 26404 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1636968456
transform 1 0 27508 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1636968456
transform 1 0 28612 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1
transform 1 0 29716 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1
transform 1 0 30268 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1636968456
transform 1 0 30452 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1636968456
transform 1 0 31556 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1636968456
transform 1 0 32660 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1636968456
transform 1 0 33764 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1
transform 1 0 34868 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1
transform 1 0 35420 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1636968456
transform 1 0 35604 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1636968456
transform 1 0 36708 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1636968456
transform 1 0 37812 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1636968456
transform 1 0 38916 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1
transform 1 0 40020 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1
transform 1 0 40572 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1636968456
transform 1 0 40756 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1636968456
transform 1 0 41860 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1636968456
transform 1 0 42964 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1636968456
transform 1 0 44068 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1
transform 1 0 45172 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1
transform 1 0 45724 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1636968456
transform 1 0 45908 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1636968456
transform 1 0 47012 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1636968456
transform 1 0 48116 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1636968456
transform 1 0 49220 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1
transform 1 0 50324 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1
transform 1 0 50876 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1636968456
transform 1 0 51060 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1636968456
transform 1 0 52164 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1636968456
transform 1 0 53268 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1636968456
transform 1 0 54372 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1
transform 1 0 55476 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1
transform 1 0 56028 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_589
timestamp 1
transform 1 0 56212 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_618
timestamp 1636968456
transform 1 0 58880 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_630
timestamp 1636968456
transform 1 0 59984 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_642
timestamp 1
transform 1 0 61088 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_645
timestamp 1636968456
transform 1 0 61364 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_657
timestamp 1636968456
transform 1 0 62468 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_669
timestamp 1636968456
transform 1 0 63572 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_681
timestamp 1636968456
transform 1 0 64676 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1
transform 1 0 65780 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1
transform 1 0 66332 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_708
timestamp 1636968456
transform 1 0 67160 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_720
timestamp 1636968456
transform 1 0 68264 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_732
timestamp 1636968456
transform 1 0 69368 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_744
timestamp 1
transform 1 0 70472 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_755
timestamp 1
transform 1 0 71484 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_757
timestamp 1636968456
transform 1 0 71668 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_769
timestamp 1636968456
transform 1 0 72772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_781
timestamp 1636968456
transform 1 0 73876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_793
timestamp 1
transform 1 0 74980 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_801
timestamp 1
transform 1 0 75716 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_807
timestamp 1
transform 1 0 76268 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_811
timestamp 1
transform 1 0 76636 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_813
timestamp 1
transform 1 0 76820 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_821
timestamp 1
transform 1 0 77556 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636968456
transform 1 0 2300 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636968456
transform 1 0 3404 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636968456
transform 1 0 4508 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1636968456
transform 1 0 5612 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1
transform 1 0 6716 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1
transform 1 0 7084 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1636968456
transform 1 0 7268 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1636968456
transform 1 0 8372 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1636968456
transform 1 0 9476 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1636968456
transform 1 0 10580 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1
transform 1 0 11684 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1
transform 1 0 12236 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1636968456
transform 1 0 12420 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1636968456
transform 1 0 13524 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1636968456
transform 1 0 14628 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1636968456
transform 1 0 15732 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1
transform 1 0 16836 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1
transform 1 0 17388 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1636968456
transform 1 0 17572 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1636968456
transform 1 0 18676 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1636968456
transform 1 0 19780 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1636968456
transform 1 0 20884 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1
transform 1 0 21988 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1
transform 1 0 22540 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1636968456
transform 1 0 22724 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1636968456
transform 1 0 23828 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1636968456
transform 1 0 24932 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1636968456
transform 1 0 26036 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1
transform 1 0 27140 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1
transform 1 0 27692 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1636968456
transform 1 0 27876 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1636968456
transform 1 0 28980 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1636968456
transform 1 0 30084 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1636968456
transform 1 0 31188 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1
transform 1 0 32292 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1
transform 1 0 32844 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1636968456
transform 1 0 33028 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1636968456
transform 1 0 34132 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1636968456
transform 1 0 35236 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1636968456
transform 1 0 36340 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1
transform 1 0 37444 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1
transform 1 0 37996 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1636968456
transform 1 0 38180 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1636968456
transform 1 0 39284 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1636968456
transform 1 0 40388 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1636968456
transform 1 0 41492 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1
transform 1 0 42596 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1
transform 1 0 43148 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1636968456
transform 1 0 43332 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1636968456
transform 1 0 44436 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1636968456
transform 1 0 45540 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1636968456
transform 1 0 46644 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1
transform 1 0 47748 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1
transform 1 0 48300 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1636968456
transform 1 0 48484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1636968456
transform 1 0 49588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1636968456
transform 1 0 50692 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1636968456
transform 1 0 51796 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1
transform 1 0 52900 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1
transform 1 0 53452 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1636968456
transform 1 0 53636 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1636968456
transform 1 0 54740 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1636968456
transform 1 0 55844 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1636968456
transform 1 0 56948 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1
transform 1 0 58052 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1
transform 1 0 58604 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_617
timestamp 1636968456
transform 1 0 58788 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_629
timestamp 1636968456
transform 1 0 59892 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_641
timestamp 1
transform 1 0 60996 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_660
timestamp 1636968456
transform 1 0 62744 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_673
timestamp 1636968456
transform 1 0 63940 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_685
timestamp 1
transform 1 0 65044 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_69_704
timestamp 1
transform 1 0 66792 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_710
timestamp 1636968456
transform 1 0 67344 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_722
timestamp 1
transform 1 0 68448 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_729
timestamp 1636968456
transform 1 0 69092 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_741
timestamp 1636968456
transform 1 0 70196 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_753
timestamp 1636968456
transform 1 0 71300 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_765
timestamp 1636968456
transform 1 0 72404 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_777
timestamp 1
transform 1 0 73508 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_783
timestamp 1
transform 1 0 74060 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_785
timestamp 1636968456
transform 1 0 74244 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_797
timestamp 1636968456
transform 1 0 75348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_809
timestamp 1636968456
transform 1 0 76452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_821
timestamp 1
transform 1 0 77556 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1636968456
transform 1 0 2300 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1636968456
transform 1 0 3404 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1
transform 1 0 4508 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636968456
transform 1 0 4692 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636968456
transform 1 0 5796 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1636968456
transform 1 0 6900 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1636968456
transform 1 0 8004 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1
transform 1 0 9108 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1
transform 1 0 9660 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1636968456
transform 1 0 9844 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1636968456
transform 1 0 10948 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1636968456
transform 1 0 12052 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1636968456
transform 1 0 13156 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1
transform 1 0 14260 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1
transform 1 0 14812 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1636968456
transform 1 0 14996 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1636968456
transform 1 0 16100 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1636968456
transform 1 0 17204 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1636968456
transform 1 0 18308 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1
transform 1 0 19412 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1
transform 1 0 19964 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1636968456
transform 1 0 20148 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1636968456
transform 1 0 21252 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1636968456
transform 1 0 22356 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1636968456
transform 1 0 23460 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1
transform 1 0 24564 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1
transform 1 0 25116 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1636968456
transform 1 0 25300 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1636968456
transform 1 0 26404 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1636968456
transform 1 0 27508 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1636968456
transform 1 0 28612 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1
transform 1 0 29716 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1
transform 1 0 30268 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1636968456
transform 1 0 30452 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1636968456
transform 1 0 31556 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1636968456
transform 1 0 32660 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1636968456
transform 1 0 33764 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1
transform 1 0 34868 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1
transform 1 0 35420 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1636968456
transform 1 0 35604 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1636968456
transform 1 0 36708 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1636968456
transform 1 0 37812 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1636968456
transform 1 0 38916 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1
transform 1 0 40020 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1
transform 1 0 40572 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1636968456
transform 1 0 40756 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1636968456
transform 1 0 41860 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1636968456
transform 1 0 42964 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1636968456
transform 1 0 44068 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1
transform 1 0 45172 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1
transform 1 0 45724 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1636968456
transform 1 0 45908 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1636968456
transform 1 0 47012 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1636968456
transform 1 0 48116 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1636968456
transform 1 0 49220 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1
transform 1 0 50324 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1
transform 1 0 50876 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1636968456
transform 1 0 51060 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1636968456
transform 1 0 52164 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1636968456
transform 1 0 53268 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1636968456
transform 1 0 54372 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1
transform 1 0 55476 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1
transform 1 0 56028 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1636968456
transform 1 0 56212 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1636968456
transform 1 0 57316 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_613
timestamp 1636968456
transform 1 0 58420 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_625
timestamp 1636968456
transform 1 0 59524 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_665
timestamp 1636968456
transform 1 0 63204 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_677
timestamp 1636968456
transform 1 0 64308 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_689
timestamp 1
transform 1 0 65412 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1
transform 1 0 66332 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_721
timestamp 1636968456
transform 1 0 68356 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_733
timestamp 1636968456
transform 1 0 69460 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_745
timestamp 1
transform 1 0 70564 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_752
timestamp 1
transform 1 0 71208 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_757
timestamp 1636968456
transform 1 0 71668 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_769
timestamp 1636968456
transform 1 0 72772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_781
timestamp 1636968456
transform 1 0 73876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_793
timestamp 1636968456
transform 1 0 74980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_805
timestamp 1
transform 1 0 76084 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_811
timestamp 1
transform 1 0 76636 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_813
timestamp 1
transform 1 0 76820 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_821
timestamp 1
transform 1 0 77556 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636968456
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636968456
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1636968456
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1636968456
transform 1 0 5612 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1
transform 1 0 6716 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1
transform 1 0 7084 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636968456
transform 1 0 7268 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1636968456
transform 1 0 8372 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1636968456
transform 1 0 9476 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1636968456
transform 1 0 10580 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1
transform 1 0 11684 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1
transform 1 0 12236 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1636968456
transform 1 0 12420 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1636968456
transform 1 0 13524 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1636968456
transform 1 0 14628 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1636968456
transform 1 0 15732 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1
transform 1 0 16836 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1
transform 1 0 17388 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1636968456
transform 1 0 17572 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1636968456
transform 1 0 18676 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1636968456
transform 1 0 19780 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1636968456
transform 1 0 20884 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1
transform 1 0 21988 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1
transform 1 0 22540 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1636968456
transform 1 0 22724 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1636968456
transform 1 0 23828 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1636968456
transform 1 0 24932 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1636968456
transform 1 0 26036 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1
transform 1 0 27140 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1
transform 1 0 27692 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1636968456
transform 1 0 27876 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1636968456
transform 1 0 28980 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1636968456
transform 1 0 30084 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1636968456
transform 1 0 31188 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1
transform 1 0 32292 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1
transform 1 0 32844 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1636968456
transform 1 0 33028 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1636968456
transform 1 0 34132 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1636968456
transform 1 0 35236 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1636968456
transform 1 0 36340 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1
transform 1 0 37444 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1
transform 1 0 37996 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1636968456
transform 1 0 38180 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1636968456
transform 1 0 39284 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1636968456
transform 1 0 40388 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1636968456
transform 1 0 41492 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1
transform 1 0 42596 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1
transform 1 0 43148 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1636968456
transform 1 0 43332 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1636968456
transform 1 0 44436 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1636968456
transform 1 0 45540 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1636968456
transform 1 0 46644 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1
transform 1 0 47748 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1
transform 1 0 48300 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1636968456
transform 1 0 48484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1636968456
transform 1 0 49588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1636968456
transform 1 0 50692 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1636968456
transform 1 0 51796 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1
transform 1 0 52900 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1
transform 1 0 53452 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1636968456
transform 1 0 53636 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1636968456
transform 1 0 54740 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1636968456
transform 1 0 55844 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1636968456
transform 1 0 56948 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1
transform 1 0 58052 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1
transform 1 0 58604 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_617
timestamp 1636968456
transform 1 0 58788 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_629
timestamp 1636968456
transform 1 0 59892 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_641
timestamp 1636968456
transform 1 0 60996 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_653
timestamp 1636968456
transform 1 0 62100 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1
transform 1 0 63204 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_671
timestamp 1
transform 1 0 63756 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_673
timestamp 1636968456
transform 1 0 63940 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_685
timestamp 1636968456
transform 1 0 65044 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_697
timestamp 1636968456
transform 1 0 66148 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_709
timestamp 1636968456
transform 1 0 67252 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_721
timestamp 1
transform 1 0 68356 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_727
timestamp 1
transform 1 0 68908 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_729
timestamp 1636968456
transform 1 0 69092 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_761
timestamp 1636968456
transform 1 0 72036 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_773
timestamp 1
transform 1 0 73140 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_781
timestamp 1
transform 1 0 73876 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_792
timestamp 1
transform 1 0 74888 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_804
timestamp 1636968456
transform 1 0 75992 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_816
timestamp 1
transform 1 0 77096 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_6
timestamp 1636968456
transform 1 0 2576 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_18
timestamp 1
transform 1 0 3680 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_26
timestamp 1
transform 1 0 4416 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636968456
transform 1 0 4692 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636968456
transform 1 0 5796 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1636968456
transform 1 0 6900 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1636968456
transform 1 0 8004 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1
transform 1 0 9108 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1
transform 1 0 9660 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1636968456
transform 1 0 9844 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1636968456
transform 1 0 10948 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1636968456
transform 1 0 12052 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1636968456
transform 1 0 13156 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1
transform 1 0 14260 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1
transform 1 0 14812 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1636968456
transform 1 0 14996 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1636968456
transform 1 0 16100 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1636968456
transform 1 0 17204 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1636968456
transform 1 0 18308 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1
transform 1 0 19412 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1
transform 1 0 19964 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1636968456
transform 1 0 20148 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1636968456
transform 1 0 21252 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1636968456
transform 1 0 22356 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1636968456
transform 1 0 23460 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1
transform 1 0 24564 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1
transform 1 0 25116 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1636968456
transform 1 0 25300 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1636968456
transform 1 0 26404 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1636968456
transform 1 0 27508 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1636968456
transform 1 0 28612 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1
transform 1 0 29716 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1
transform 1 0 30268 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1636968456
transform 1 0 30452 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1636968456
transform 1 0 31556 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1636968456
transform 1 0 32660 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1636968456
transform 1 0 33764 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1
transform 1 0 34868 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1
transform 1 0 35420 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1636968456
transform 1 0 35604 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1636968456
transform 1 0 36708 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1636968456
transform 1 0 37812 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1636968456
transform 1 0 38916 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1
transform 1 0 40020 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1
transform 1 0 40572 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1636968456
transform 1 0 40756 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1636968456
transform 1 0 41860 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1636968456
transform 1 0 42964 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1636968456
transform 1 0 44068 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1
transform 1 0 45172 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1
transform 1 0 45724 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1636968456
transform 1 0 45908 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1636968456
transform 1 0 47012 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1636968456
transform 1 0 48116 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1636968456
transform 1 0 49220 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1
transform 1 0 50324 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1
transform 1 0 50876 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1636968456
transform 1 0 51060 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1636968456
transform 1 0 52164 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1636968456
transform 1 0 53268 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1636968456
transform 1 0 54372 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1
transform 1 0 55476 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1
transform 1 0 56028 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1636968456
transform 1 0 56212 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1636968456
transform 1 0 57316 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1636968456
transform 1 0 58420 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_625
timestamp 1636968456
transform 1 0 59524 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_637
timestamp 1
transform 1 0 60628 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1
transform 1 0 61180 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_645
timestamp 1636968456
transform 1 0 61364 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_657
timestamp 1636968456
transform 1 0 62468 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_669
timestamp 1
transform 1 0 63572 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_677
timestamp 1
transform 1 0 64308 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_683
timestamp 1636968456
transform 1 0 64860 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_695
timestamp 1
transform 1 0 65964 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1
transform 1 0 66332 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_701
timestamp 1636968456
transform 1 0 66516 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_713
timestamp 1636968456
transform 1 0 67620 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_725
timestamp 1636968456
transform 1 0 68724 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_737
timestamp 1636968456
transform 1 0 69828 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_749
timestamp 1
transform 1 0 70932 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_754
timestamp 1
transform 1 0 71392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_757
timestamp 1636968456
transform 1 0 71668 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_769
timestamp 1636968456
transform 1 0 72772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_781
timestamp 1
transform 1 0 73876 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_785
timestamp 1
transform 1 0 74244 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_809
timestamp 1
transform 1 0 76452 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_813
timestamp 1
transform 1 0 76820 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_821
timestamp 1
transform 1 0 77556 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636968456
transform 1 0 2300 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636968456
transform 1 0 3404 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636968456
transform 1 0 4508 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1636968456
transform 1 0 5612 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1
transform 1 0 6716 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1
transform 1 0 7084 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1636968456
transform 1 0 7268 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1636968456
transform 1 0 8372 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1636968456
transform 1 0 9476 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1636968456
transform 1 0 10580 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1
transform 1 0 11684 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1
transform 1 0 12236 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1636968456
transform 1 0 12420 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1636968456
transform 1 0 13524 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1636968456
transform 1 0 14628 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1636968456
transform 1 0 15732 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1
transform 1 0 16836 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1
transform 1 0 17388 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1636968456
transform 1 0 17572 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1636968456
transform 1 0 18676 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1636968456
transform 1 0 19780 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1636968456
transform 1 0 20884 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1
transform 1 0 21988 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1
transform 1 0 22540 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1636968456
transform 1 0 22724 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1636968456
transform 1 0 23828 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1636968456
transform 1 0 24932 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1636968456
transform 1 0 26036 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1
transform 1 0 27140 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1
transform 1 0 27692 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1636968456
transform 1 0 27876 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1636968456
transform 1 0 28980 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1636968456
transform 1 0 30084 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1636968456
transform 1 0 31188 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1
transform 1 0 32292 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1
transform 1 0 32844 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1636968456
transform 1 0 33028 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1636968456
transform 1 0 34132 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1636968456
transform 1 0 35236 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1636968456
transform 1 0 36340 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1
transform 1 0 37444 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1
transform 1 0 37996 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1636968456
transform 1 0 38180 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1636968456
transform 1 0 39284 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1636968456
transform 1 0 40388 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1636968456
transform 1 0 41492 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1
transform 1 0 42596 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1
transform 1 0 43148 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1636968456
transform 1 0 43332 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1636968456
transform 1 0 44436 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1636968456
transform 1 0 45540 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1636968456
transform 1 0 46644 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1
transform 1 0 47748 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1
transform 1 0 48300 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1636968456
transform 1 0 48484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1636968456
transform 1 0 49588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1636968456
transform 1 0 50692 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1636968456
transform 1 0 51796 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1
transform 1 0 52900 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1
transform 1 0 53452 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1636968456
transform 1 0 53636 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1636968456
transform 1 0 54740 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1636968456
transform 1 0 55844 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_597
timestamp 1
transform 1 0 56948 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_605
timestamp 1
transform 1 0 57684 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_611
timestamp 1
transform 1 0 58236 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1
transform 1 0 58604 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_620
timestamp 1636968456
transform 1 0 59064 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_632
timestamp 1636968456
transform 1 0 60168 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_644
timestamp 1636968456
transform 1 0 61272 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_656
timestamp 1636968456
transform 1 0 62376 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_668
timestamp 1
transform 1 0 63480 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_673
timestamp 1636968456
transform 1 0 63940 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_685
timestamp 1636968456
transform 1 0 65044 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_697
timestamp 1636968456
transform 1 0 66148 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_709
timestamp 1636968456
transform 1 0 67252 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_721
timestamp 1
transform 1 0 68356 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_727
timestamp 1
transform 1 0 68908 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_729
timestamp 1636968456
transform 1 0 69092 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_741
timestamp 1636968456
transform 1 0 70196 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_753
timestamp 1636968456
transform 1 0 71300 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_765
timestamp 1636968456
transform 1 0 72404 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_777
timestamp 1
transform 1 0 73508 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_783
timestamp 1
transform 1 0 74060 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_785
timestamp 1636968456
transform 1 0 74244 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_797
timestamp 1636968456
transform 1 0 75348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_809
timestamp 1636968456
transform 1 0 76452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_821
timestamp 1
transform 1 0 77556 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636968456
transform 1 0 2300 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636968456
transform 1 0 3404 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1
transform 1 0 4508 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636968456
transform 1 0 4692 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1636968456
transform 1 0 5796 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1636968456
transform 1 0 6900 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1636968456
transform 1 0 8004 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1
transform 1 0 9108 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1
transform 1 0 9660 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1636968456
transform 1 0 9844 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1636968456
transform 1 0 10948 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1636968456
transform 1 0 12052 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1636968456
transform 1 0 13156 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1
transform 1 0 14260 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1
transform 1 0 14812 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1636968456
transform 1 0 14996 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1636968456
transform 1 0 16100 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1636968456
transform 1 0 17204 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1636968456
transform 1 0 18308 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1
transform 1 0 19412 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1
transform 1 0 19964 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1636968456
transform 1 0 20148 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1636968456
transform 1 0 21252 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1636968456
transform 1 0 22356 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1636968456
transform 1 0 23460 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1
transform 1 0 24564 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1
transform 1 0 25116 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1636968456
transform 1 0 25300 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1636968456
transform 1 0 26404 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1636968456
transform 1 0 27508 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1636968456
transform 1 0 28612 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1
transform 1 0 29716 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1
transform 1 0 30268 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1636968456
transform 1 0 30452 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1636968456
transform 1 0 31556 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1636968456
transform 1 0 32660 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1636968456
transform 1 0 33764 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1
transform 1 0 34868 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1
transform 1 0 35420 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1636968456
transform 1 0 35604 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1636968456
transform 1 0 36708 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1636968456
transform 1 0 37812 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1636968456
transform 1 0 38916 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1
transform 1 0 40020 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1
transform 1 0 40572 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1636968456
transform 1 0 40756 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1636968456
transform 1 0 41860 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1636968456
transform 1 0 42964 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1636968456
transform 1 0 44068 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1
transform 1 0 45172 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1
transform 1 0 45724 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1636968456
transform 1 0 45908 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1636968456
transform 1 0 47012 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1636968456
transform 1 0 48116 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1636968456
transform 1 0 49220 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1
transform 1 0 50324 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1
transform 1 0 50876 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1636968456
transform 1 0 51060 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1636968456
transform 1 0 52164 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1636968456
transform 1 0 53268 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1636968456
transform 1 0 54372 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1
transform 1 0 55476 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1
transform 1 0 56028 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1636968456
transform 1 0 56212 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_601
timestamp 1
transform 1 0 57316 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_633
timestamp 1
transform 1 0 60260 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_641
timestamp 1
transform 1 0 60996 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_645
timestamp 1636968456
transform 1 0 61364 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_657
timestamp 1636968456
transform 1 0 62468 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_669
timestamp 1636968456
transform 1 0 63572 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_681
timestamp 1636968456
transform 1 0 64676 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1
transform 1 0 65780 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1
transform 1 0 66332 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_701
timestamp 1636968456
transform 1 0 66516 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_713
timestamp 1636968456
transform 1 0 67620 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_725
timestamp 1636968456
transform 1 0 68724 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_737
timestamp 1636968456
transform 1 0 69828 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_749
timestamp 1
transform 1 0 70932 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_755
timestamp 1
transform 1 0 71484 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_757
timestamp 1636968456
transform 1 0 71668 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_769
timestamp 1636968456
transform 1 0 72772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_781
timestamp 1636968456
transform 1 0 73876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_793
timestamp 1636968456
transform 1 0 74980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_805
timestamp 1
transform 1 0 76084 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_811
timestamp 1
transform 1 0 76636 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_813
timestamp 1
transform 1 0 76820 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_821
timestamp 1
transform 1 0 77556 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636968456
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636968456
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1636968456
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1636968456
transform 1 0 5612 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1
transform 1 0 6716 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1
transform 1 0 7084 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1636968456
transform 1 0 7268 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1636968456
transform 1 0 8372 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1636968456
transform 1 0 9476 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1636968456
transform 1 0 10580 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1
transform 1 0 11684 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1
transform 1 0 12236 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1636968456
transform 1 0 12420 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1636968456
transform 1 0 13524 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1636968456
transform 1 0 14628 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1636968456
transform 1 0 15732 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1
transform 1 0 16836 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1
transform 1 0 17388 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1636968456
transform 1 0 17572 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1636968456
transform 1 0 18676 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1636968456
transform 1 0 19780 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1636968456
transform 1 0 20884 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1
transform 1 0 21988 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1
transform 1 0 22540 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1636968456
transform 1 0 22724 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1636968456
transform 1 0 23828 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1636968456
transform 1 0 24932 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1636968456
transform 1 0 26036 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1
transform 1 0 27140 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1
transform 1 0 27692 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1636968456
transform 1 0 27876 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1636968456
transform 1 0 28980 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1636968456
transform 1 0 30084 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1636968456
transform 1 0 31188 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1
transform 1 0 32292 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1
transform 1 0 32844 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1636968456
transform 1 0 33028 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1636968456
transform 1 0 34132 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1636968456
transform 1 0 35236 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1636968456
transform 1 0 36340 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1
transform 1 0 37444 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1
transform 1 0 37996 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1636968456
transform 1 0 38180 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1636968456
transform 1 0 39284 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1636968456
transform 1 0 40388 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1636968456
transform 1 0 41492 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1
transform 1 0 42596 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1
transform 1 0 43148 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1636968456
transform 1 0 43332 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1636968456
transform 1 0 44436 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1636968456
transform 1 0 45540 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1636968456
transform 1 0 46644 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1
transform 1 0 47748 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1
transform 1 0 48300 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1636968456
transform 1 0 48484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1636968456
transform 1 0 49588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1636968456
transform 1 0 50692 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1636968456
transform 1 0 51796 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1
transform 1 0 52900 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1
transform 1 0 53452 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1636968456
transform 1 0 53636 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1636968456
transform 1 0 54740 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1636968456
transform 1 0 55844 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1636968456
transform 1 0 56948 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1
transform 1 0 58052 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1
transform 1 0 58604 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_617
timestamp 1636968456
transform 1 0 58788 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_629
timestamp 1636968456
transform 1 0 59892 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_641
timestamp 1636968456
transform 1 0 60996 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_653
timestamp 1636968456
transform 1 0 62100 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1
transform 1 0 63204 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1
transform 1 0 63756 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_673
timestamp 1636968456
transform 1 0 63940 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_685
timestamp 1
transform 1 0 65044 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_709
timestamp 1636968456
transform 1 0 67252 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_721
timestamp 1
transform 1 0 68356 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_727
timestamp 1
transform 1 0 68908 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_729
timestamp 1636968456
transform 1 0 69092 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_741
timestamp 1636968456
transform 1 0 70196 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_753
timestamp 1636968456
transform 1 0 71300 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_765
timestamp 1636968456
transform 1 0 72404 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_777
timestamp 1
transform 1 0 73508 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_783
timestamp 1
transform 1 0 74060 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_785
timestamp 1636968456
transform 1 0 74244 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_797
timestamp 1636968456
transform 1 0 75348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_809
timestamp 1636968456
transform 1 0 76452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_821
timestamp 1
transform 1 0 77556 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636968456
transform 1 0 2300 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636968456
transform 1 0 3404 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1
transform 1 0 4508 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1636968456
transform 1 0 4692 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1636968456
transform 1 0 5796 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1636968456
transform 1 0 6900 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1636968456
transform 1 0 8004 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1
transform 1 0 9108 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1
transform 1 0 9660 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1636968456
transform 1 0 9844 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1636968456
transform 1 0 10948 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1636968456
transform 1 0 12052 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1636968456
transform 1 0 13156 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1
transform 1 0 14260 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1
transform 1 0 14812 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1636968456
transform 1 0 14996 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1636968456
transform 1 0 16100 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1636968456
transform 1 0 17204 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1636968456
transform 1 0 18308 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1
transform 1 0 19412 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1
transform 1 0 19964 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1636968456
transform 1 0 20148 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1636968456
transform 1 0 21252 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1636968456
transform 1 0 22356 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1636968456
transform 1 0 23460 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1
transform 1 0 24564 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1
transform 1 0 25116 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1636968456
transform 1 0 25300 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1636968456
transform 1 0 26404 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1636968456
transform 1 0 27508 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1636968456
transform 1 0 28612 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1
transform 1 0 29716 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1
transform 1 0 30268 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1636968456
transform 1 0 30452 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1636968456
transform 1 0 31556 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1636968456
transform 1 0 32660 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1636968456
transform 1 0 33764 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1
transform 1 0 34868 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1
transform 1 0 35420 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1636968456
transform 1 0 35604 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1636968456
transform 1 0 36708 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1636968456
transform 1 0 37812 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1636968456
transform 1 0 38916 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1
transform 1 0 40020 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1
transform 1 0 40572 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1636968456
transform 1 0 40756 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1636968456
transform 1 0 41860 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1636968456
transform 1 0 42964 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1636968456
transform 1 0 44068 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1
transform 1 0 45172 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1
transform 1 0 45724 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1636968456
transform 1 0 45908 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1636968456
transform 1 0 47012 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1636968456
transform 1 0 48116 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1636968456
transform 1 0 49220 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1
transform 1 0 50324 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1
transform 1 0 50876 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1636968456
transform 1 0 51060 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1636968456
transform 1 0 52164 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1636968456
transform 1 0 53268 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1636968456
transform 1 0 54372 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1
transform 1 0 55476 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1
transform 1 0 56028 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1636968456
transform 1 0 56212 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1636968456
transform 1 0 57316 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1636968456
transform 1 0 58420 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_625
timestamp 1636968456
transform 1 0 59524 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1
transform 1 0 60628 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1
transform 1 0 61180 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_645
timestamp 1636968456
transform 1 0 61364 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_657
timestamp 1636968456
transform 1 0 62468 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_669
timestamp 1636968456
transform 1 0 63572 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_681
timestamp 1
transform 1 0 64676 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_689
timestamp 1
transform 1 0 65412 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_697
timestamp 1
transform 1 0 66148 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_709
timestamp 1636968456
transform 1 0 67252 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_721
timestamp 1636968456
transform 1 0 68356 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_733
timestamp 1636968456
transform 1 0 69460 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_745
timestamp 1
transform 1 0 70564 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_753
timestamp 1
transform 1 0 71300 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_757
timestamp 1636968456
transform 1 0 71668 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_769
timestamp 1636968456
transform 1 0 72772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_781
timestamp 1636968456
transform 1 0 73876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_793
timestamp 1636968456
transform 1 0 74980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_805
timestamp 1
transform 1 0 76084 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_811
timestamp 1
transform 1 0 76636 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_813
timestamp 1
transform 1 0 76820 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_821
timestamp 1
transform 1 0 77556 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1636968456
transform 1 0 2300 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1636968456
transform 1 0 3404 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1636968456
transform 1 0 4508 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1636968456
transform 1 0 5612 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1
transform 1 0 6716 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1
transform 1 0 7084 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1636968456
transform 1 0 7268 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1636968456
transform 1 0 8372 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1636968456
transform 1 0 9476 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1636968456
transform 1 0 10580 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1
transform 1 0 11684 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1
transform 1 0 12236 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1636968456
transform 1 0 12420 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1636968456
transform 1 0 13524 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1636968456
transform 1 0 14628 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1636968456
transform 1 0 15732 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1
transform 1 0 16836 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1
transform 1 0 17388 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1636968456
transform 1 0 17572 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1636968456
transform 1 0 18676 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1636968456
transform 1 0 19780 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1636968456
transform 1 0 20884 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1
transform 1 0 21988 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1
transform 1 0 22540 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1636968456
transform 1 0 22724 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1636968456
transform 1 0 23828 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1636968456
transform 1 0 24932 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1636968456
transform 1 0 26036 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1
transform 1 0 27140 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1
transform 1 0 27692 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1636968456
transform 1 0 27876 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1636968456
transform 1 0 28980 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1636968456
transform 1 0 30084 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1636968456
transform 1 0 31188 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1
transform 1 0 32292 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1
transform 1 0 32844 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1636968456
transform 1 0 33028 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1636968456
transform 1 0 34132 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1636968456
transform 1 0 35236 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1636968456
transform 1 0 36340 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1
transform 1 0 37444 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1
transform 1 0 37996 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1636968456
transform 1 0 38180 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1636968456
transform 1 0 39284 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1636968456
transform 1 0 40388 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1636968456
transform 1 0 41492 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1
transform 1 0 42596 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1
transform 1 0 43148 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1636968456
transform 1 0 43332 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1636968456
transform 1 0 44436 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1636968456
transform 1 0 45540 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1636968456
transform 1 0 46644 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1
transform 1 0 47748 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1
transform 1 0 48300 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1636968456
transform 1 0 48484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1636968456
transform 1 0 49588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1636968456
transform 1 0 50692 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1636968456
transform 1 0 51796 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1
transform 1 0 52900 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1
transform 1 0 53452 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1636968456
transform 1 0 53636 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1636968456
transform 1 0 54740 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1636968456
transform 1 0 55844 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1636968456
transform 1 0 56948 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1
transform 1 0 58052 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1
transform 1 0 58604 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_617
timestamp 1636968456
transform 1 0 58788 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_629
timestamp 1636968456
transform 1 0 59892 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_641
timestamp 1636968456
transform 1 0 60996 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_653
timestamp 1636968456
transform 1 0 62100 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1
transform 1 0 63204 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1
transform 1 0 63756 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_673
timestamp 1636968456
transform 1 0 63940 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_685
timestamp 1636968456
transform 1 0 65044 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_697
timestamp 1636968456
transform 1 0 66148 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_709
timestamp 1636968456
transform 1 0 67252 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_721
timestamp 1
transform 1 0 68356 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_727
timestamp 1
transform 1 0 68908 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_729
timestamp 1636968456
transform 1 0 69092 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_741
timestamp 1636968456
transform 1 0 70196 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_753
timestamp 1636968456
transform 1 0 71300 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_765
timestamp 1636968456
transform 1 0 72404 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_777
timestamp 1
transform 1 0 73508 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_783
timestamp 1
transform 1 0 74060 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_785
timestamp 1636968456
transform 1 0 74244 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_797
timestamp 1636968456
transform 1 0 75348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_809
timestamp 1636968456
transform 1 0 76452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_821
timestamp 1
transform 1 0 77556 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636968456
transform 1 0 2300 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636968456
transform 1 0 3404 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1
transform 1 0 4508 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1636968456
transform 1 0 4692 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1636968456
transform 1 0 5796 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1636968456
transform 1 0 6900 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1636968456
transform 1 0 8004 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1
transform 1 0 9108 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1
transform 1 0 9660 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1636968456
transform 1 0 9844 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1636968456
transform 1 0 10948 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1636968456
transform 1 0 12052 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1636968456
transform 1 0 13156 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1
transform 1 0 14260 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1
transform 1 0 14812 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1636968456
transform 1 0 14996 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1636968456
transform 1 0 16100 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1636968456
transform 1 0 17204 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1636968456
transform 1 0 18308 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1
transform 1 0 19412 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1
transform 1 0 19964 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1636968456
transform 1 0 20148 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1636968456
transform 1 0 21252 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1636968456
transform 1 0 22356 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1636968456
transform 1 0 23460 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1
transform 1 0 24564 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1
transform 1 0 25116 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1636968456
transform 1 0 25300 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1636968456
transform 1 0 26404 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1636968456
transform 1 0 27508 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1636968456
transform 1 0 28612 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1
transform 1 0 29716 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1
transform 1 0 30268 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1636968456
transform 1 0 30452 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1636968456
transform 1 0 31556 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1636968456
transform 1 0 32660 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1636968456
transform 1 0 33764 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1
transform 1 0 34868 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1
transform 1 0 35420 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1636968456
transform 1 0 35604 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1636968456
transform 1 0 36708 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1636968456
transform 1 0 37812 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1636968456
transform 1 0 38916 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1
transform 1 0 40020 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1
transform 1 0 40572 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1636968456
transform 1 0 40756 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1636968456
transform 1 0 41860 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1636968456
transform 1 0 42964 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1636968456
transform 1 0 44068 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1
transform 1 0 45172 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1
transform 1 0 45724 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1636968456
transform 1 0 45908 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1636968456
transform 1 0 47012 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1636968456
transform 1 0 48116 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1636968456
transform 1 0 49220 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1
transform 1 0 50324 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1
transform 1 0 50876 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1636968456
transform 1 0 51060 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1636968456
transform 1 0 52164 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1636968456
transform 1 0 53268 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1636968456
transform 1 0 54372 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1
transform 1 0 55476 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1
transform 1 0 56028 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1636968456
transform 1 0 56212 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1636968456
transform 1 0 57316 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1636968456
transform 1 0 58420 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_625
timestamp 1636968456
transform 1 0 59524 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1
transform 1 0 60628 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1
transform 1 0 61180 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_645
timestamp 1636968456
transform 1 0 61364 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_657
timestamp 1636968456
transform 1 0 62468 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_669
timestamp 1636968456
transform 1 0 63572 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_681
timestamp 1636968456
transform 1 0 64676 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1
transform 1 0 65780 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1
transform 1 0 66332 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_701
timestamp 1636968456
transform 1 0 66516 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_713
timestamp 1636968456
transform 1 0 67620 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_725
timestamp 1636968456
transform 1 0 68724 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_737
timestamp 1636968456
transform 1 0 69828 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_749
timestamp 1
transform 1 0 70932 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_755
timestamp 1
transform 1 0 71484 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_757
timestamp 1636968456
transform 1 0 71668 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_769
timestamp 1636968456
transform 1 0 72772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_781
timestamp 1636968456
transform 1 0 73876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_793
timestamp 1636968456
transform 1 0 74980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_805
timestamp 1
transform 1 0 76084 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_811
timestamp 1
transform 1 0 76636 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_813
timestamp 1
transform 1 0 76820 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_821
timestamp 1
transform 1 0 77556 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636968456
transform 1 0 2300 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636968456
transform 1 0 3404 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1636968456
transform 1 0 4508 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1636968456
transform 1 0 5612 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1
transform 1 0 6716 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1
transform 1 0 7084 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1636968456
transform 1 0 7268 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1636968456
transform 1 0 8372 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1636968456
transform 1 0 9476 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1636968456
transform 1 0 10580 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1
transform 1 0 11684 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1
transform 1 0 12236 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1636968456
transform 1 0 12420 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1636968456
transform 1 0 13524 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1636968456
transform 1 0 14628 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1636968456
transform 1 0 15732 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1
transform 1 0 16836 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1
transform 1 0 17388 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1636968456
transform 1 0 17572 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1636968456
transform 1 0 18676 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1636968456
transform 1 0 19780 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1636968456
transform 1 0 20884 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1
transform 1 0 21988 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1
transform 1 0 22540 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1636968456
transform 1 0 22724 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1636968456
transform 1 0 23828 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1636968456
transform 1 0 24932 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1636968456
transform 1 0 26036 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1
transform 1 0 27140 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1
transform 1 0 27692 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1636968456
transform 1 0 27876 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1636968456
transform 1 0 28980 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1636968456
transform 1 0 30084 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1636968456
transform 1 0 31188 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1
transform 1 0 32292 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1
transform 1 0 32844 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1636968456
transform 1 0 33028 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1636968456
transform 1 0 34132 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1636968456
transform 1 0 35236 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1636968456
transform 1 0 36340 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1
transform 1 0 37444 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1
transform 1 0 37996 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1636968456
transform 1 0 38180 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1636968456
transform 1 0 39284 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1636968456
transform 1 0 40388 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1636968456
transform 1 0 41492 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1
transform 1 0 42596 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1
transform 1 0 43148 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1636968456
transform 1 0 43332 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1636968456
transform 1 0 44436 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1636968456
transform 1 0 45540 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1636968456
transform 1 0 46644 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1
transform 1 0 47748 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1
transform 1 0 48300 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1636968456
transform 1 0 48484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1636968456
transform 1 0 49588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1636968456
transform 1 0 50692 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1636968456
transform 1 0 51796 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1
transform 1 0 52900 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1
transform 1 0 53452 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1636968456
transform 1 0 53636 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1636968456
transform 1 0 54740 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1636968456
transform 1 0 55844 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1636968456
transform 1 0 56948 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1
transform 1 0 58052 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1
transform 1 0 58604 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_617
timestamp 1636968456
transform 1 0 58788 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_629
timestamp 1636968456
transform 1 0 59892 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_641
timestamp 1636968456
transform 1 0 60996 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_653
timestamp 1636968456
transform 1 0 62100 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1
transform 1 0 63204 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1
transform 1 0 63756 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_673
timestamp 1636968456
transform 1 0 63940 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_685
timestamp 1636968456
transform 1 0 65044 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_697
timestamp 1636968456
transform 1 0 66148 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_709
timestamp 1636968456
transform 1 0 67252 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_721
timestamp 1
transform 1 0 68356 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_727
timestamp 1
transform 1 0 68908 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_729
timestamp 1636968456
transform 1 0 69092 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_741
timestamp 1636968456
transform 1 0 70196 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_753
timestamp 1636968456
transform 1 0 71300 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_765
timestamp 1636968456
transform 1 0 72404 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_777
timestamp 1
transform 1 0 73508 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_783
timestamp 1
transform 1 0 74060 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_785
timestamp 1636968456
transform 1 0 74244 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_797
timestamp 1636968456
transform 1 0 75348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_809
timestamp 1636968456
transform 1 0 76452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_821
timestamp 1
transform 1 0 77556 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636968456
transform 1 0 2300 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636968456
transform 1 0 3404 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1
transform 1 0 4508 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1636968456
transform 1 0 4692 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1636968456
transform 1 0 5796 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1636968456
transform 1 0 6900 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1636968456
transform 1 0 8004 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1
transform 1 0 9108 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1
transform 1 0 9660 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1636968456
transform 1 0 9844 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1636968456
transform 1 0 10948 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1636968456
transform 1 0 12052 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1636968456
transform 1 0 13156 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1
transform 1 0 14260 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1
transform 1 0 14812 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1636968456
transform 1 0 14996 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1636968456
transform 1 0 16100 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1636968456
transform 1 0 17204 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1636968456
transform 1 0 18308 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1
transform 1 0 19412 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1
transform 1 0 19964 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1636968456
transform 1 0 20148 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1636968456
transform 1 0 21252 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1636968456
transform 1 0 22356 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1636968456
transform 1 0 23460 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1
transform 1 0 24564 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1
transform 1 0 25116 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1636968456
transform 1 0 25300 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1636968456
transform 1 0 26404 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1636968456
transform 1 0 27508 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1636968456
transform 1 0 28612 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1
transform 1 0 29716 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1
transform 1 0 30268 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1636968456
transform 1 0 30452 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1636968456
transform 1 0 31556 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1636968456
transform 1 0 32660 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1636968456
transform 1 0 33764 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1
transform 1 0 34868 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1
transform 1 0 35420 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1636968456
transform 1 0 35604 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1636968456
transform 1 0 36708 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1636968456
transform 1 0 37812 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1636968456
transform 1 0 38916 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1
transform 1 0 40020 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1
transform 1 0 40572 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1636968456
transform 1 0 40756 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1636968456
transform 1 0 41860 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1636968456
transform 1 0 42964 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1636968456
transform 1 0 44068 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1
transform 1 0 45172 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1
transform 1 0 45724 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1636968456
transform 1 0 45908 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1636968456
transform 1 0 47012 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1636968456
transform 1 0 48116 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1636968456
transform 1 0 49220 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1
transform 1 0 50324 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1
transform 1 0 50876 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1636968456
transform 1 0 51060 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1636968456
transform 1 0 52164 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1636968456
transform 1 0 53268 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1636968456
transform 1 0 54372 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1
transform 1 0 55476 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1
transform 1 0 56028 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1636968456
transform 1 0 56212 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1636968456
transform 1 0 57316 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1636968456
transform 1 0 58420 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_625
timestamp 1636968456
transform 1 0 59524 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1
transform 1 0 60628 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1
transform 1 0 61180 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_645
timestamp 1636968456
transform 1 0 61364 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_657
timestamp 1636968456
transform 1 0 62468 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_669
timestamp 1636968456
transform 1 0 63572 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_681
timestamp 1636968456
transform 1 0 64676 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_693
timestamp 1
transform 1 0 65780 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_699
timestamp 1
transform 1 0 66332 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_701
timestamp 1636968456
transform 1 0 66516 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_713
timestamp 1636968456
transform 1 0 67620 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_725
timestamp 1636968456
transform 1 0 68724 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_737
timestamp 1636968456
transform 1 0 69828 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_749
timestamp 1
transform 1 0 70932 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_755
timestamp 1
transform 1 0 71484 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_757
timestamp 1636968456
transform 1 0 71668 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_769
timestamp 1636968456
transform 1 0 72772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_781
timestamp 1636968456
transform 1 0 73876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_793
timestamp 1636968456
transform 1 0 74980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_805
timestamp 1
transform 1 0 76084 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_811
timestamp 1
transform 1 0 76636 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_813
timestamp 1
transform 1 0 76820 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_821
timestamp 1
transform 1 0 77556 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636968456
transform 1 0 2300 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636968456
transform 1 0 3404 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1636968456
transform 1 0 4508 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1636968456
transform 1 0 5612 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1
transform 1 0 6716 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1
transform 1 0 7084 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1636968456
transform 1 0 7268 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1636968456
transform 1 0 8372 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1636968456
transform 1 0 9476 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1636968456
transform 1 0 10580 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1
transform 1 0 11684 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1
transform 1 0 12236 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1636968456
transform 1 0 12420 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1636968456
transform 1 0 13524 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1636968456
transform 1 0 14628 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1636968456
transform 1 0 15732 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1
transform 1 0 16836 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1
transform 1 0 17388 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1636968456
transform 1 0 17572 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1636968456
transform 1 0 18676 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1636968456
transform 1 0 19780 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1636968456
transform 1 0 20884 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1
transform 1 0 21988 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1
transform 1 0 22540 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1636968456
transform 1 0 22724 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1636968456
transform 1 0 23828 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1636968456
transform 1 0 24932 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1636968456
transform 1 0 26036 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1
transform 1 0 27140 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1
transform 1 0 27692 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1636968456
transform 1 0 27876 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1636968456
transform 1 0 28980 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1636968456
transform 1 0 30084 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1636968456
transform 1 0 31188 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1
transform 1 0 32292 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1
transform 1 0 32844 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1636968456
transform 1 0 33028 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1636968456
transform 1 0 34132 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1636968456
transform 1 0 35236 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1636968456
transform 1 0 36340 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1
transform 1 0 37444 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1
transform 1 0 37996 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1636968456
transform 1 0 38180 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1636968456
transform 1 0 39284 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1636968456
transform 1 0 40388 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1636968456
transform 1 0 41492 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1
transform 1 0 42596 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1
transform 1 0 43148 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1636968456
transform 1 0 43332 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1636968456
transform 1 0 44436 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1636968456
transform 1 0 45540 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1636968456
transform 1 0 46644 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1
transform 1 0 47748 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1
transform 1 0 48300 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1636968456
transform 1 0 48484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1636968456
transform 1 0 49588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1636968456
transform 1 0 50692 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1636968456
transform 1 0 51796 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1
transform 1 0 52900 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1
transform 1 0 53452 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1636968456
transform 1 0 53636 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1636968456
transform 1 0 54740 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1636968456
transform 1 0 55844 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1636968456
transform 1 0 56948 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1
transform 1 0 58052 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1
transform 1 0 58604 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_617
timestamp 1636968456
transform 1 0 58788 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_629
timestamp 1636968456
transform 1 0 59892 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_641
timestamp 1636968456
transform 1 0 60996 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_653
timestamp 1636968456
transform 1 0 62100 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_665
timestamp 1
transform 1 0 63204 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_671
timestamp 1
transform 1 0 63756 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_673
timestamp 1636968456
transform 1 0 63940 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_685
timestamp 1636968456
transform 1 0 65044 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_697
timestamp 1636968456
transform 1 0 66148 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_709
timestamp 1636968456
transform 1 0 67252 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_721
timestamp 1
transform 1 0 68356 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_727
timestamp 1
transform 1 0 68908 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_729
timestamp 1636968456
transform 1 0 69092 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_741
timestamp 1636968456
transform 1 0 70196 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_753
timestamp 1636968456
transform 1 0 71300 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_765
timestamp 1636968456
transform 1 0 72404 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_777
timestamp 1
transform 1 0 73508 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_783
timestamp 1
transform 1 0 74060 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_785
timestamp 1636968456
transform 1 0 74244 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_797
timestamp 1636968456
transform 1 0 75348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_809
timestamp 1636968456
transform 1 0 76452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_821
timestamp 1
transform 1 0 77556 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1636968456
transform 1 0 2300 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1636968456
transform 1 0 3404 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1
transform 1 0 4508 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1636968456
transform 1 0 4692 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1636968456
transform 1 0 5796 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1636968456
transform 1 0 6900 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1636968456
transform 1 0 8004 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1
transform 1 0 9108 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1
transform 1 0 9660 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1636968456
transform 1 0 9844 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1636968456
transform 1 0 10948 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1636968456
transform 1 0 12052 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1636968456
transform 1 0 13156 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1
transform 1 0 14260 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1
transform 1 0 14812 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1636968456
transform 1 0 14996 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1636968456
transform 1 0 16100 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1636968456
transform 1 0 17204 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1636968456
transform 1 0 18308 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1
transform 1 0 19412 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1
transform 1 0 19964 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1636968456
transform 1 0 20148 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1636968456
transform 1 0 21252 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1636968456
transform 1 0 22356 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1636968456
transform 1 0 23460 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1
transform 1 0 24564 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1
transform 1 0 25116 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1636968456
transform 1 0 25300 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1636968456
transform 1 0 26404 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1636968456
transform 1 0 27508 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1636968456
transform 1 0 28612 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1
transform 1 0 29716 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1
transform 1 0 30268 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1636968456
transform 1 0 30452 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1636968456
transform 1 0 31556 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1636968456
transform 1 0 32660 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1636968456
transform 1 0 33764 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1
transform 1 0 34868 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1
transform 1 0 35420 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1636968456
transform 1 0 35604 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1636968456
transform 1 0 36708 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1636968456
transform 1 0 37812 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1636968456
transform 1 0 38916 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1
transform 1 0 40020 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1
transform 1 0 40572 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1636968456
transform 1 0 40756 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1636968456
transform 1 0 41860 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1636968456
transform 1 0 42964 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1636968456
transform 1 0 44068 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1
transform 1 0 45172 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1
transform 1 0 45724 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1636968456
transform 1 0 45908 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1636968456
transform 1 0 47012 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1636968456
transform 1 0 48116 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1636968456
transform 1 0 49220 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1
transform 1 0 50324 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1
transform 1 0 50876 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1636968456
transform 1 0 51060 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1636968456
transform 1 0 52164 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1636968456
transform 1 0 53268 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1636968456
transform 1 0 54372 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1
transform 1 0 55476 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1
transform 1 0 56028 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1636968456
transform 1 0 56212 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1636968456
transform 1 0 57316 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1636968456
transform 1 0 58420 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_625
timestamp 1636968456
transform 1 0 59524 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_637
timestamp 1
transform 1 0 60628 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_643
timestamp 1
transform 1 0 61180 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_645
timestamp 1636968456
transform 1 0 61364 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_657
timestamp 1636968456
transform 1 0 62468 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_669
timestamp 1636968456
transform 1 0 63572 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_681
timestamp 1636968456
transform 1 0 64676 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_693
timestamp 1
transform 1 0 65780 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_699
timestamp 1
transform 1 0 66332 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_701
timestamp 1636968456
transform 1 0 66516 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_713
timestamp 1636968456
transform 1 0 67620 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_725
timestamp 1636968456
transform 1 0 68724 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_737
timestamp 1636968456
transform 1 0 69828 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_749
timestamp 1
transform 1 0 70932 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_755
timestamp 1
transform 1 0 71484 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_757
timestamp 1636968456
transform 1 0 71668 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_769
timestamp 1636968456
transform 1 0 72772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_781
timestamp 1636968456
transform 1 0 73876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_793
timestamp 1636968456
transform 1 0 74980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_805
timestamp 1
transform 1 0 76084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_811
timestamp 1
transform 1 0 76636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_813
timestamp 1
transform 1 0 76820 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_821
timestamp 1
transform 1 0 77556 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636968456
transform 1 0 2300 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636968456
transform 1 0 3404 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1636968456
transform 1 0 4508 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1636968456
transform 1 0 5612 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1
transform 1 0 6716 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1
transform 1 0 7084 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1636968456
transform 1 0 7268 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1636968456
transform 1 0 8372 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1636968456
transform 1 0 9476 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1636968456
transform 1 0 10580 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1
transform 1 0 11684 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1
transform 1 0 12236 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1636968456
transform 1 0 12420 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1636968456
transform 1 0 13524 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1636968456
transform 1 0 14628 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1636968456
transform 1 0 15732 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1
transform 1 0 16836 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1
transform 1 0 17388 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1636968456
transform 1 0 17572 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1636968456
transform 1 0 18676 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1636968456
transform 1 0 19780 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1636968456
transform 1 0 20884 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1
transform 1 0 21988 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1
transform 1 0 22540 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1636968456
transform 1 0 22724 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1636968456
transform 1 0 23828 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1636968456
transform 1 0 24932 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1636968456
transform 1 0 26036 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1
transform 1 0 27140 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1
transform 1 0 27692 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1636968456
transform 1 0 27876 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1636968456
transform 1 0 28980 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1636968456
transform 1 0 30084 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1636968456
transform 1 0 31188 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1
transform 1 0 32292 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1
transform 1 0 32844 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1636968456
transform 1 0 33028 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1636968456
transform 1 0 34132 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1636968456
transform 1 0 35236 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1636968456
transform 1 0 36340 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1
transform 1 0 37444 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1
transform 1 0 37996 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1636968456
transform 1 0 38180 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1636968456
transform 1 0 39284 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1636968456
transform 1 0 40388 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1636968456
transform 1 0 41492 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1
transform 1 0 42596 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1
transform 1 0 43148 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1636968456
transform 1 0 43332 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1636968456
transform 1 0 44436 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1636968456
transform 1 0 45540 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1636968456
transform 1 0 46644 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1
transform 1 0 47748 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1
transform 1 0 48300 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1636968456
transform 1 0 48484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1636968456
transform 1 0 49588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1636968456
transform 1 0 50692 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1636968456
transform 1 0 51796 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1
transform 1 0 52900 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1
transform 1 0 53452 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1636968456
transform 1 0 53636 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1636968456
transform 1 0 54740 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1636968456
transform 1 0 55844 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1636968456
transform 1 0 56948 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1
transform 1 0 58052 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1
transform 1 0 58604 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_617
timestamp 1636968456
transform 1 0 58788 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_629
timestamp 1636968456
transform 1 0 59892 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_641
timestamp 1636968456
transform 1 0 60996 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_653
timestamp 1636968456
transform 1 0 62100 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_665
timestamp 1
transform 1 0 63204 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_671
timestamp 1
transform 1 0 63756 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_673
timestamp 1636968456
transform 1 0 63940 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_685
timestamp 1636968456
transform 1 0 65044 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_697
timestamp 1636968456
transform 1 0 66148 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_709
timestamp 1636968456
transform 1 0 67252 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_721
timestamp 1
transform 1 0 68356 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_727
timestamp 1
transform 1 0 68908 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_729
timestamp 1636968456
transform 1 0 69092 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_741
timestamp 1636968456
transform 1 0 70196 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_753
timestamp 1636968456
transform 1 0 71300 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_765
timestamp 1636968456
transform 1 0 72404 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_777
timestamp 1
transform 1 0 73508 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_783
timestamp 1
transform 1 0 74060 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_785
timestamp 1636968456
transform 1 0 74244 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_797
timestamp 1636968456
transform 1 0 75348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_809
timestamp 1636968456
transform 1 0 76452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_821
timestamp 1
transform 1 0 77556 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636968456
transform 1 0 2300 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636968456
transform 1 0 3404 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1
transform 1 0 4508 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1636968456
transform 1 0 4692 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1636968456
transform 1 0 5796 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1636968456
transform 1 0 6900 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1636968456
transform 1 0 8004 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1
transform 1 0 9108 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1
transform 1 0 9660 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1636968456
transform 1 0 9844 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1636968456
transform 1 0 10948 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1636968456
transform 1 0 12052 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1636968456
transform 1 0 13156 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1
transform 1 0 14260 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1
transform 1 0 14812 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1636968456
transform 1 0 14996 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1636968456
transform 1 0 16100 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1636968456
transform 1 0 17204 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1636968456
transform 1 0 18308 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1
transform 1 0 19412 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1
transform 1 0 19964 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1636968456
transform 1 0 20148 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1636968456
transform 1 0 21252 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1636968456
transform 1 0 22356 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1636968456
transform 1 0 23460 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1
transform 1 0 24564 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1
transform 1 0 25116 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1636968456
transform 1 0 25300 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1636968456
transform 1 0 26404 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1636968456
transform 1 0 27508 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1636968456
transform 1 0 28612 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1
transform 1 0 29716 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1
transform 1 0 30268 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1636968456
transform 1 0 30452 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1636968456
transform 1 0 31556 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1636968456
transform 1 0 32660 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1636968456
transform 1 0 33764 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1
transform 1 0 34868 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1
transform 1 0 35420 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1636968456
transform 1 0 35604 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1636968456
transform 1 0 36708 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1636968456
transform 1 0 37812 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1636968456
transform 1 0 38916 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1
transform 1 0 40020 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1
transform 1 0 40572 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1636968456
transform 1 0 40756 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1636968456
transform 1 0 41860 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1636968456
transform 1 0 42964 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1636968456
transform 1 0 44068 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1
transform 1 0 45172 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1
transform 1 0 45724 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1636968456
transform 1 0 45908 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1636968456
transform 1 0 47012 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1636968456
transform 1 0 48116 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1636968456
transform 1 0 49220 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1
transform 1 0 50324 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1
transform 1 0 50876 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1636968456
transform 1 0 51060 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1636968456
transform 1 0 52164 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1636968456
transform 1 0 53268 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1636968456
transform 1 0 54372 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1
transform 1 0 55476 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1
transform 1 0 56028 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1636968456
transform 1 0 56212 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1636968456
transform 1 0 57316 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1636968456
transform 1 0 58420 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_625
timestamp 1636968456
transform 1 0 59524 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1
transform 1 0 60628 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1
transform 1 0 61180 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_645
timestamp 1636968456
transform 1 0 61364 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_657
timestamp 1636968456
transform 1 0 62468 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_669
timestamp 1636968456
transform 1 0 63572 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_681
timestamp 1636968456
transform 1 0 64676 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1
transform 1 0 65780 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1
transform 1 0 66332 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_701
timestamp 1636968456
transform 1 0 66516 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_713
timestamp 1636968456
transform 1 0 67620 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_725
timestamp 1636968456
transform 1 0 68724 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_737
timestamp 1636968456
transform 1 0 69828 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_749
timestamp 1
transform 1 0 70932 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_755
timestamp 1
transform 1 0 71484 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_757
timestamp 1636968456
transform 1 0 71668 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_769
timestamp 1636968456
transform 1 0 72772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_781
timestamp 1636968456
transform 1 0 73876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_793
timestamp 1636968456
transform 1 0 74980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_805
timestamp 1
transform 1 0 76084 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_811
timestamp 1
transform 1 0 76636 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_813
timestamp 1
transform 1 0 76820 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_821
timestamp 1
transform 1 0 77556 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1636968456
transform 1 0 2300 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1636968456
transform 1 0 3404 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1636968456
transform 1 0 4508 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1636968456
transform 1 0 5612 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1
transform 1 0 6716 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1
transform 1 0 7084 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1636968456
transform 1 0 7268 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1636968456
transform 1 0 8372 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1636968456
transform 1 0 9476 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1636968456
transform 1 0 10580 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1
transform 1 0 11684 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1
transform 1 0 12236 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1636968456
transform 1 0 12420 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1636968456
transform 1 0 13524 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1636968456
transform 1 0 14628 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1636968456
transform 1 0 15732 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1
transform 1 0 16836 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1
transform 1 0 17388 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1636968456
transform 1 0 17572 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1636968456
transform 1 0 18676 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1636968456
transform 1 0 19780 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1636968456
transform 1 0 20884 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1
transform 1 0 21988 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1
transform 1 0 22540 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1636968456
transform 1 0 22724 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1636968456
transform 1 0 23828 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1636968456
transform 1 0 24932 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1636968456
transform 1 0 26036 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1
transform 1 0 27140 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1
transform 1 0 27692 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1636968456
transform 1 0 27876 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1636968456
transform 1 0 28980 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1636968456
transform 1 0 30084 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1636968456
transform 1 0 31188 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1
transform 1 0 32292 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1
transform 1 0 32844 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1636968456
transform 1 0 33028 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1636968456
transform 1 0 34132 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1636968456
transform 1 0 35236 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1636968456
transform 1 0 36340 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1
transform 1 0 37444 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1
transform 1 0 37996 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1636968456
transform 1 0 38180 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1636968456
transform 1 0 39284 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1636968456
transform 1 0 40388 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1636968456
transform 1 0 41492 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1
transform 1 0 42596 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1
transform 1 0 43148 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1636968456
transform 1 0 43332 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1636968456
transform 1 0 44436 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1636968456
transform 1 0 45540 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1636968456
transform 1 0 46644 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1
transform 1 0 47748 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1
transform 1 0 48300 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1636968456
transform 1 0 48484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1636968456
transform 1 0 49588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1636968456
transform 1 0 50692 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1636968456
transform 1 0 51796 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1
transform 1 0 52900 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1
transform 1 0 53452 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1636968456
transform 1 0 53636 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1636968456
transform 1 0 54740 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1636968456
transform 1 0 55844 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1636968456
transform 1 0 56948 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1
transform 1 0 58052 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1
transform 1 0 58604 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_617
timestamp 1636968456
transform 1 0 58788 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_629
timestamp 1636968456
transform 1 0 59892 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_641
timestamp 1636968456
transform 1 0 60996 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_653
timestamp 1636968456
transform 1 0 62100 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1
transform 1 0 63204 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1
transform 1 0 63756 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_673
timestamp 1636968456
transform 1 0 63940 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_685
timestamp 1636968456
transform 1 0 65044 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_697
timestamp 1636968456
transform 1 0 66148 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_709
timestamp 1636968456
transform 1 0 67252 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_721
timestamp 1
transform 1 0 68356 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_727
timestamp 1
transform 1 0 68908 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_729
timestamp 1636968456
transform 1 0 69092 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_741
timestamp 1636968456
transform 1 0 70196 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_753
timestamp 1636968456
transform 1 0 71300 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_765
timestamp 1636968456
transform 1 0 72404 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_777
timestamp 1
transform 1 0 73508 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_783
timestamp 1
transform 1 0 74060 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_785
timestamp 1636968456
transform 1 0 74244 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_797
timestamp 1636968456
transform 1 0 75348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_809
timestamp 1636968456
transform 1 0 76452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_821
timestamp 1
transform 1 0 77556 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636968456
transform 1 0 2300 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636968456
transform 1 0 3404 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1
transform 1 0 4508 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1636968456
transform 1 0 4692 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1636968456
transform 1 0 5796 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1636968456
transform 1 0 6900 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1636968456
transform 1 0 8004 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1
transform 1 0 9108 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1
transform 1 0 9660 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1636968456
transform 1 0 9844 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1636968456
transform 1 0 10948 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1636968456
transform 1 0 12052 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1636968456
transform 1 0 13156 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1
transform 1 0 14260 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1
transform 1 0 14812 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1636968456
transform 1 0 14996 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1636968456
transform 1 0 16100 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1636968456
transform 1 0 17204 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1636968456
transform 1 0 18308 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1
transform 1 0 19412 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1
transform 1 0 19964 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1636968456
transform 1 0 20148 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1636968456
transform 1 0 21252 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1636968456
transform 1 0 22356 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1636968456
transform 1 0 23460 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1
transform 1 0 24564 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1
transform 1 0 25116 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1636968456
transform 1 0 25300 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1636968456
transform 1 0 26404 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1636968456
transform 1 0 27508 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1636968456
transform 1 0 28612 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1
transform 1 0 29716 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1
transform 1 0 30268 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1636968456
transform 1 0 30452 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1636968456
transform 1 0 31556 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1636968456
transform 1 0 32660 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1636968456
transform 1 0 33764 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1
transform 1 0 34868 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1
transform 1 0 35420 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1636968456
transform 1 0 35604 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1636968456
transform 1 0 36708 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1636968456
transform 1 0 37812 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1636968456
transform 1 0 38916 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1
transform 1 0 40020 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1
transform 1 0 40572 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1636968456
transform 1 0 40756 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1636968456
transform 1 0 41860 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1636968456
transform 1 0 42964 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1636968456
transform 1 0 44068 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1
transform 1 0 45172 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1
transform 1 0 45724 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1636968456
transform 1 0 45908 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1636968456
transform 1 0 47012 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1636968456
transform 1 0 48116 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1636968456
transform 1 0 49220 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1
transform 1 0 50324 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1
transform 1 0 50876 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1636968456
transform 1 0 51060 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1636968456
transform 1 0 52164 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1636968456
transform 1 0 53268 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1636968456
transform 1 0 54372 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1
transform 1 0 55476 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1
transform 1 0 56028 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1636968456
transform 1 0 56212 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1636968456
transform 1 0 57316 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1636968456
transform 1 0 58420 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_625
timestamp 1636968456
transform 1 0 59524 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1
transform 1 0 60628 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1
transform 1 0 61180 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_645
timestamp 1636968456
transform 1 0 61364 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_657
timestamp 1636968456
transform 1 0 62468 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_669
timestamp 1636968456
transform 1 0 63572 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_681
timestamp 1636968456
transform 1 0 64676 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1
transform 1 0 65780 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1
transform 1 0 66332 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_701
timestamp 1636968456
transform 1 0 66516 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_713
timestamp 1636968456
transform 1 0 67620 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_725
timestamp 1636968456
transform 1 0 68724 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_737
timestamp 1636968456
transform 1 0 69828 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_749
timestamp 1
transform 1 0 70932 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_755
timestamp 1
transform 1 0 71484 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_757
timestamp 1636968456
transform 1 0 71668 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_769
timestamp 1636968456
transform 1 0 72772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_781
timestamp 1636968456
transform 1 0 73876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_793
timestamp 1636968456
transform 1 0 74980 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_805
timestamp 1
transform 1 0 76084 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_811
timestamp 1
transform 1 0 76636 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_813
timestamp 1
transform 1 0 76820 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_821
timestamp 1
transform 1 0 77556 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1636968456
transform 1 0 2300 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1636968456
transform 1 0 3404 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1636968456
transform 1 0 4508 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1636968456
transform 1 0 5612 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1
transform 1 0 6716 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1
transform 1 0 7084 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1636968456
transform 1 0 7268 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1636968456
transform 1 0 8372 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1636968456
transform 1 0 9476 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1636968456
transform 1 0 10580 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1
transform 1 0 11684 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1
transform 1 0 12236 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1636968456
transform 1 0 12420 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1636968456
transform 1 0 13524 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1636968456
transform 1 0 14628 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1636968456
transform 1 0 15732 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1
transform 1 0 16836 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1
transform 1 0 17388 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1636968456
transform 1 0 17572 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1636968456
transform 1 0 18676 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1636968456
transform 1 0 19780 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1636968456
transform 1 0 20884 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1
transform 1 0 21988 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1
transform 1 0 22540 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1636968456
transform 1 0 22724 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1636968456
transform 1 0 23828 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1636968456
transform 1 0 24932 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1636968456
transform 1 0 26036 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1
transform 1 0 27140 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1
transform 1 0 27692 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1636968456
transform 1 0 27876 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1636968456
transform 1 0 28980 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1636968456
transform 1 0 30084 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1636968456
transform 1 0 31188 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1
transform 1 0 32292 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1
transform 1 0 32844 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1636968456
transform 1 0 33028 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1636968456
transform 1 0 34132 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1636968456
transform 1 0 35236 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1636968456
transform 1 0 36340 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1
transform 1 0 37444 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1
transform 1 0 37996 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1636968456
transform 1 0 38180 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1636968456
transform 1 0 39284 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1636968456
transform 1 0 40388 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1636968456
transform 1 0 41492 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1
transform 1 0 42596 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1
transform 1 0 43148 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1636968456
transform 1 0 43332 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1636968456
transform 1 0 44436 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1636968456
transform 1 0 45540 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1636968456
transform 1 0 46644 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1
transform 1 0 47748 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1
transform 1 0 48300 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1636968456
transform 1 0 48484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1636968456
transform 1 0 49588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1636968456
transform 1 0 50692 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1636968456
transform 1 0 51796 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1
transform 1 0 52900 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1
transform 1 0 53452 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1636968456
transform 1 0 53636 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1636968456
transform 1 0 54740 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1636968456
transform 1 0 55844 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1636968456
transform 1 0 56948 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1
transform 1 0 58052 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1
transform 1 0 58604 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_617
timestamp 1636968456
transform 1 0 58788 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_629
timestamp 1636968456
transform 1 0 59892 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_641
timestamp 1636968456
transform 1 0 60996 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_653
timestamp 1636968456
transform 1 0 62100 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1
transform 1 0 63204 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1
transform 1 0 63756 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_673
timestamp 1636968456
transform 1 0 63940 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_685
timestamp 1636968456
transform 1 0 65044 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_697
timestamp 1636968456
transform 1 0 66148 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_709
timestamp 1636968456
transform 1 0 67252 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_721
timestamp 1
transform 1 0 68356 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_727
timestamp 1
transform 1 0 68908 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_729
timestamp 1636968456
transform 1 0 69092 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_741
timestamp 1636968456
transform 1 0 70196 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_753
timestamp 1636968456
transform 1 0 71300 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_765
timestamp 1636968456
transform 1 0 72404 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_777
timestamp 1
transform 1 0 73508 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_783
timestamp 1
transform 1 0 74060 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_785
timestamp 1636968456
transform 1 0 74244 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_797
timestamp 1636968456
transform 1 0 75348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_809
timestamp 1
transform 1 0 76452 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_817
timestamp 1
transform 1 0 77188 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1636968456
transform 1 0 2300 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1636968456
transform 1 0 3404 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1
transform 1 0 4508 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1636968456
transform 1 0 4692 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1636968456
transform 1 0 5796 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1636968456
transform 1 0 6900 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1636968456
transform 1 0 8004 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1
transform 1 0 9108 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1
transform 1 0 9660 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1636968456
transform 1 0 9844 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1636968456
transform 1 0 10948 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1636968456
transform 1 0 12052 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1636968456
transform 1 0 13156 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1
transform 1 0 14260 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1
transform 1 0 14812 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1636968456
transform 1 0 14996 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1636968456
transform 1 0 16100 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1636968456
transform 1 0 17204 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1636968456
transform 1 0 18308 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1
transform 1 0 19412 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1
transform 1 0 19964 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1636968456
transform 1 0 20148 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1636968456
transform 1 0 21252 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1636968456
transform 1 0 22356 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1636968456
transform 1 0 23460 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1
transform 1 0 24564 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1
transform 1 0 25116 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1636968456
transform 1 0 25300 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1636968456
transform 1 0 26404 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1636968456
transform 1 0 27508 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1636968456
transform 1 0 28612 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1
transform 1 0 29716 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1
transform 1 0 30268 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1636968456
transform 1 0 30452 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1636968456
transform 1 0 31556 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1636968456
transform 1 0 32660 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1636968456
transform 1 0 33764 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1
transform 1 0 34868 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1
transform 1 0 35420 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1636968456
transform 1 0 35604 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1636968456
transform 1 0 36708 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1636968456
transform 1 0 37812 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1636968456
transform 1 0 38916 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1
transform 1 0 40020 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1
transform 1 0 40572 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1636968456
transform 1 0 40756 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1636968456
transform 1 0 41860 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1636968456
transform 1 0 42964 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1636968456
transform 1 0 44068 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1
transform 1 0 45172 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1
transform 1 0 45724 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1636968456
transform 1 0 45908 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1636968456
transform 1 0 47012 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1636968456
transform 1 0 48116 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1636968456
transform 1 0 49220 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1
transform 1 0 50324 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1
transform 1 0 50876 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1636968456
transform 1 0 51060 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1636968456
transform 1 0 52164 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1636968456
transform 1 0 53268 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1636968456
transform 1 0 54372 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1
transform 1 0 55476 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1
transform 1 0 56028 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1636968456
transform 1 0 56212 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1636968456
transform 1 0 57316 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1636968456
transform 1 0 58420 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_625
timestamp 1636968456
transform 1 0 59524 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1
transform 1 0 60628 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1
transform 1 0 61180 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_645
timestamp 1636968456
transform 1 0 61364 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_657
timestamp 1636968456
transform 1 0 62468 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_669
timestamp 1636968456
transform 1 0 63572 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_681
timestamp 1636968456
transform 1 0 64676 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_693
timestamp 1
transform 1 0 65780 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_699
timestamp 1
transform 1 0 66332 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_701
timestamp 1636968456
transform 1 0 66516 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_713
timestamp 1636968456
transform 1 0 67620 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_725
timestamp 1636968456
transform 1 0 68724 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_737
timestamp 1636968456
transform 1 0 69828 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_749
timestamp 1
transform 1 0 70932 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_755
timestamp 1
transform 1 0 71484 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_757
timestamp 1636968456
transform 1 0 71668 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_769
timestamp 1636968456
transform 1 0 72772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_781
timestamp 1636968456
transform 1 0 73876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_793
timestamp 1636968456
transform 1 0 74980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_805
timestamp 1
transform 1 0 76084 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_811
timestamp 1
transform 1 0 76636 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_813
timestamp 1
transform 1 0 76820 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_821
timestamp 1
transform 1 0 77556 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1636968456
transform 1 0 2300 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1636968456
transform 1 0 3404 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1636968456
transform 1 0 4508 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1636968456
transform 1 0 5612 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1
transform 1 0 6716 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1
transform 1 0 7084 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1636968456
transform 1 0 7268 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1636968456
transform 1 0 8372 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1636968456
transform 1 0 9476 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1636968456
transform 1 0 10580 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1
transform 1 0 11684 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1
transform 1 0 12236 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1636968456
transform 1 0 12420 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1636968456
transform 1 0 13524 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1636968456
transform 1 0 14628 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1636968456
transform 1 0 15732 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1
transform 1 0 16836 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1
transform 1 0 17388 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1636968456
transform 1 0 17572 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1636968456
transform 1 0 18676 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1636968456
transform 1 0 19780 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1636968456
transform 1 0 20884 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1
transform 1 0 21988 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1
transform 1 0 22540 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1636968456
transform 1 0 22724 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1636968456
transform 1 0 23828 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1636968456
transform 1 0 24932 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1636968456
transform 1 0 26036 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1
transform 1 0 27140 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1
transform 1 0 27692 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1636968456
transform 1 0 27876 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1636968456
transform 1 0 28980 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1636968456
transform 1 0 30084 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1636968456
transform 1 0 31188 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1
transform 1 0 32292 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1
transform 1 0 32844 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1636968456
transform 1 0 33028 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1636968456
transform 1 0 34132 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1636968456
transform 1 0 35236 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1636968456
transform 1 0 36340 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1
transform 1 0 37444 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1
transform 1 0 37996 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1636968456
transform 1 0 38180 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1636968456
transform 1 0 39284 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1636968456
transform 1 0 40388 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1636968456
transform 1 0 41492 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1
transform 1 0 42596 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1
transform 1 0 43148 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1636968456
transform 1 0 43332 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1636968456
transform 1 0 44436 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1636968456
transform 1 0 45540 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1636968456
transform 1 0 46644 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1
transform 1 0 47748 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1
transform 1 0 48300 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1636968456
transform 1 0 48484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1636968456
transform 1 0 49588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1636968456
transform 1 0 50692 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1636968456
transform 1 0 51796 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1
transform 1 0 52900 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1
transform 1 0 53452 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1636968456
transform 1 0 53636 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1636968456
transform 1 0 54740 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1636968456
transform 1 0 55844 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1636968456
transform 1 0 56948 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1
transform 1 0 58052 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1
transform 1 0 58604 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_617
timestamp 1636968456
transform 1 0 58788 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_629
timestamp 1636968456
transform 1 0 59892 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_641
timestamp 1636968456
transform 1 0 60996 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_653
timestamp 1636968456
transform 1 0 62100 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1
transform 1 0 63204 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1
transform 1 0 63756 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_673
timestamp 1636968456
transform 1 0 63940 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_685
timestamp 1636968456
transform 1 0 65044 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_697
timestamp 1636968456
transform 1 0 66148 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_709
timestamp 1636968456
transform 1 0 67252 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_721
timestamp 1
transform 1 0 68356 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_727
timestamp 1
transform 1 0 68908 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_729
timestamp 1636968456
transform 1 0 69092 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_741
timestamp 1636968456
transform 1 0 70196 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_753
timestamp 1636968456
transform 1 0 71300 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_765
timestamp 1636968456
transform 1 0 72404 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_777
timestamp 1
transform 1 0 73508 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_783
timestamp 1
transform 1 0 74060 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_785
timestamp 1636968456
transform 1 0 74244 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_797
timestamp 1636968456
transform 1 0 75348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_809
timestamp 1636968456
transform 1 0 76452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_821
timestamp 1
transform 1 0 77556 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1636968456
transform 1 0 2300 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1636968456
transform 1 0 3404 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1
transform 1 0 4508 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1636968456
transform 1 0 4692 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1636968456
transform 1 0 5796 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1636968456
transform 1 0 6900 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1636968456
transform 1 0 8004 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1
transform 1 0 9108 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1
transform 1 0 9660 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1636968456
transform 1 0 9844 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1636968456
transform 1 0 10948 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1636968456
transform 1 0 12052 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1636968456
transform 1 0 13156 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1
transform 1 0 14260 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1
transform 1 0 14812 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1636968456
transform 1 0 14996 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1636968456
transform 1 0 16100 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1636968456
transform 1 0 17204 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1636968456
transform 1 0 18308 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1
transform 1 0 19412 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1
transform 1 0 19964 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1636968456
transform 1 0 20148 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1636968456
transform 1 0 21252 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1636968456
transform 1 0 22356 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1636968456
transform 1 0 23460 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1
transform 1 0 24564 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1
transform 1 0 25116 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1636968456
transform 1 0 25300 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1636968456
transform 1 0 26404 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1636968456
transform 1 0 27508 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1636968456
transform 1 0 28612 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1
transform 1 0 29716 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1
transform 1 0 30268 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1636968456
transform 1 0 30452 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1636968456
transform 1 0 31556 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1636968456
transform 1 0 32660 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1636968456
transform 1 0 33764 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1
transform 1 0 34868 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1
transform 1 0 35420 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1636968456
transform 1 0 35604 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1636968456
transform 1 0 36708 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1636968456
transform 1 0 37812 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1636968456
transform 1 0 38916 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1
transform 1 0 40020 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1
transform 1 0 40572 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1636968456
transform 1 0 40756 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1636968456
transform 1 0 41860 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1636968456
transform 1 0 42964 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1636968456
transform 1 0 44068 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1
transform 1 0 45172 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1
transform 1 0 45724 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1636968456
transform 1 0 45908 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1636968456
transform 1 0 47012 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1636968456
transform 1 0 48116 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1636968456
transform 1 0 49220 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1
transform 1 0 50324 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1
transform 1 0 50876 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1636968456
transform 1 0 51060 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1636968456
transform 1 0 52164 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1636968456
transform 1 0 53268 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1636968456
transform 1 0 54372 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1
transform 1 0 55476 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1
transform 1 0 56028 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1636968456
transform 1 0 56212 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1636968456
transform 1 0 57316 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1636968456
transform 1 0 58420 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_625
timestamp 1636968456
transform 1 0 59524 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1
transform 1 0 60628 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1
transform 1 0 61180 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_645
timestamp 1636968456
transform 1 0 61364 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_657
timestamp 1636968456
transform 1 0 62468 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_669
timestamp 1636968456
transform 1 0 63572 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_681
timestamp 1636968456
transform 1 0 64676 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1
transform 1 0 65780 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1
transform 1 0 66332 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_701
timestamp 1636968456
transform 1 0 66516 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_713
timestamp 1636968456
transform 1 0 67620 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_725
timestamp 1636968456
transform 1 0 68724 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_737
timestamp 1636968456
transform 1 0 69828 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_749
timestamp 1
transform 1 0 70932 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_755
timestamp 1
transform 1 0 71484 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_757
timestamp 1636968456
transform 1 0 71668 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_769
timestamp 1636968456
transform 1 0 72772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_781
timestamp 1636968456
transform 1 0 73876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_793
timestamp 1636968456
transform 1 0 74980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_805
timestamp 1
transform 1 0 76084 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_811
timestamp 1
transform 1 0 76636 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_813
timestamp 1
transform 1 0 76820 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_821
timestamp 1
transform 1 0 77556 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1636968456
transform 1 0 2300 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1636968456
transform 1 0 3404 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1636968456
transform 1 0 4508 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1636968456
transform 1 0 5612 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1
transform 1 0 6716 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1
transform 1 0 7084 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1636968456
transform 1 0 7268 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1636968456
transform 1 0 8372 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1636968456
transform 1 0 9476 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1636968456
transform 1 0 10580 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1
transform 1 0 11684 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1
transform 1 0 12236 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1636968456
transform 1 0 12420 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1636968456
transform 1 0 13524 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1636968456
transform 1 0 14628 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1636968456
transform 1 0 15732 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1
transform 1 0 16836 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1
transform 1 0 17388 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1636968456
transform 1 0 17572 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1636968456
transform 1 0 18676 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1636968456
transform 1 0 19780 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1636968456
transform 1 0 20884 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1
transform 1 0 21988 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1
transform 1 0 22540 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1636968456
transform 1 0 22724 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1636968456
transform 1 0 23828 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1636968456
transform 1 0 24932 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1636968456
transform 1 0 26036 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1
transform 1 0 27140 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1
transform 1 0 27692 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1636968456
transform 1 0 27876 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1636968456
transform 1 0 28980 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1636968456
transform 1 0 30084 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1636968456
transform 1 0 31188 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1
transform 1 0 32292 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1
transform 1 0 32844 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1636968456
transform 1 0 33028 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1636968456
transform 1 0 34132 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1636968456
transform 1 0 35236 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1636968456
transform 1 0 36340 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1
transform 1 0 37444 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1
transform 1 0 37996 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1636968456
transform 1 0 38180 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1636968456
transform 1 0 39284 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1636968456
transform 1 0 40388 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1636968456
transform 1 0 41492 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1
transform 1 0 42596 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1
transform 1 0 43148 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1636968456
transform 1 0 43332 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1636968456
transform 1 0 44436 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1636968456
transform 1 0 45540 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1636968456
transform 1 0 46644 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1
transform 1 0 47748 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1
transform 1 0 48300 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1636968456
transform 1 0 48484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1636968456
transform 1 0 49588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1636968456
transform 1 0 50692 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1636968456
transform 1 0 51796 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1
transform 1 0 52900 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1
transform 1 0 53452 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1636968456
transform 1 0 53636 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1636968456
transform 1 0 54740 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1636968456
transform 1 0 55844 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1636968456
transform 1 0 56948 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1
transform 1 0 58052 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1
transform 1 0 58604 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_617
timestamp 1636968456
transform 1 0 58788 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_629
timestamp 1636968456
transform 1 0 59892 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_641
timestamp 1636968456
transform 1 0 60996 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_653
timestamp 1636968456
transform 1 0 62100 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1
transform 1 0 63204 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1
transform 1 0 63756 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_673
timestamp 1636968456
transform 1 0 63940 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_685
timestamp 1636968456
transform 1 0 65044 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_697
timestamp 1636968456
transform 1 0 66148 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_709
timestamp 1636968456
transform 1 0 67252 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_721
timestamp 1
transform 1 0 68356 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_727
timestamp 1
transform 1 0 68908 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_729
timestamp 1636968456
transform 1 0 69092 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_741
timestamp 1636968456
transform 1 0 70196 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_753
timestamp 1636968456
transform 1 0 71300 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_765
timestamp 1636968456
transform 1 0 72404 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_777
timestamp 1
transform 1 0 73508 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_783
timestamp 1
transform 1 0 74060 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_785
timestamp 1636968456
transform 1 0 74244 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_797
timestamp 1636968456
transform 1 0 75348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_809
timestamp 1
transform 1 0 76452 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_817
timestamp 1
transform 1 0 77188 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1636968456
transform 1 0 2300 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1636968456
transform 1 0 3404 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1
transform 1 0 4508 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1636968456
transform 1 0 4692 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1636968456
transform 1 0 5796 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1636968456
transform 1 0 6900 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1636968456
transform 1 0 8004 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1
transform 1 0 9108 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1
transform 1 0 9660 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1636968456
transform 1 0 9844 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1636968456
transform 1 0 10948 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1636968456
transform 1 0 12052 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1636968456
transform 1 0 13156 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1
transform 1 0 14260 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1
transform 1 0 14812 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1636968456
transform 1 0 14996 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1636968456
transform 1 0 16100 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1636968456
transform 1 0 17204 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1636968456
transform 1 0 18308 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1
transform 1 0 19412 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1
transform 1 0 19964 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1636968456
transform 1 0 20148 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1636968456
transform 1 0 21252 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1636968456
transform 1 0 22356 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1636968456
transform 1 0 23460 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1
transform 1 0 24564 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1
transform 1 0 25116 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1636968456
transform 1 0 25300 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1636968456
transform 1 0 26404 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1636968456
transform 1 0 27508 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1636968456
transform 1 0 28612 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1
transform 1 0 29716 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1
transform 1 0 30268 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1636968456
transform 1 0 30452 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1636968456
transform 1 0 31556 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1636968456
transform 1 0 32660 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1636968456
transform 1 0 33764 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1
transform 1 0 34868 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1
transform 1 0 35420 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1636968456
transform 1 0 35604 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1636968456
transform 1 0 36708 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1636968456
transform 1 0 37812 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1636968456
transform 1 0 38916 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1
transform 1 0 40020 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1
transform 1 0 40572 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1636968456
transform 1 0 40756 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1636968456
transform 1 0 41860 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1636968456
transform 1 0 42964 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1636968456
transform 1 0 44068 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1
transform 1 0 45172 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1
transform 1 0 45724 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1636968456
transform 1 0 45908 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1636968456
transform 1 0 47012 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1636968456
transform 1 0 48116 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1636968456
transform 1 0 49220 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1
transform 1 0 50324 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1
transform 1 0 50876 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1636968456
transform 1 0 51060 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1636968456
transform 1 0 52164 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1636968456
transform 1 0 53268 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1636968456
transform 1 0 54372 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1
transform 1 0 55476 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1
transform 1 0 56028 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1636968456
transform 1 0 56212 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1636968456
transform 1 0 57316 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1636968456
transform 1 0 58420 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_625
timestamp 1636968456
transform 1 0 59524 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1
transform 1 0 60628 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1
transform 1 0 61180 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_645
timestamp 1636968456
transform 1 0 61364 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_657
timestamp 1636968456
transform 1 0 62468 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_669
timestamp 1636968456
transform 1 0 63572 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_681
timestamp 1636968456
transform 1 0 64676 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1
transform 1 0 65780 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1
transform 1 0 66332 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_701
timestamp 1636968456
transform 1 0 66516 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_713
timestamp 1636968456
transform 1 0 67620 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_725
timestamp 1636968456
transform 1 0 68724 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_737
timestamp 1636968456
transform 1 0 69828 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_749
timestamp 1
transform 1 0 70932 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_755
timestamp 1
transform 1 0 71484 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_757
timestamp 1636968456
transform 1 0 71668 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_769
timestamp 1636968456
transform 1 0 72772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_781
timestamp 1636968456
transform 1 0 73876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_793
timestamp 1636968456
transform 1 0 74980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_805
timestamp 1
transform 1 0 76084 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_811
timestamp 1
transform 1 0 76636 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_813
timestamp 1
transform 1 0 76820 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_821
timestamp 1
transform 1 0 77556 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1636968456
transform 1 0 2300 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1636968456
transform 1 0 3404 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1636968456
transform 1 0 4508 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1636968456
transform 1 0 5612 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1
transform 1 0 6716 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1
transform 1 0 7084 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1636968456
transform 1 0 7268 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1636968456
transform 1 0 8372 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1636968456
transform 1 0 9476 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1636968456
transform 1 0 10580 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1
transform 1 0 11684 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1
transform 1 0 12236 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1636968456
transform 1 0 12420 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1636968456
transform 1 0 13524 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1636968456
transform 1 0 14628 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1636968456
transform 1 0 15732 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1
transform 1 0 16836 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1
transform 1 0 17388 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1636968456
transform 1 0 17572 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1636968456
transform 1 0 18676 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1636968456
transform 1 0 19780 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1636968456
transform 1 0 20884 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1
transform 1 0 21988 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1
transform 1 0 22540 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1636968456
transform 1 0 22724 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1636968456
transform 1 0 23828 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1636968456
transform 1 0 24932 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1636968456
transform 1 0 26036 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1
transform 1 0 27140 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1
transform 1 0 27692 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1636968456
transform 1 0 27876 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1636968456
transform 1 0 28980 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1636968456
transform 1 0 30084 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1636968456
transform 1 0 31188 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1
transform 1 0 32292 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1
transform 1 0 32844 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1636968456
transform 1 0 33028 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1636968456
transform 1 0 34132 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1636968456
transform 1 0 35236 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1636968456
transform 1 0 36340 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1
transform 1 0 37444 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1
transform 1 0 37996 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1636968456
transform 1 0 38180 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1636968456
transform 1 0 39284 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1636968456
transform 1 0 40388 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1636968456
transform 1 0 41492 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1
transform 1 0 42596 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1
transform 1 0 43148 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1636968456
transform 1 0 43332 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1636968456
transform 1 0 44436 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1636968456
transform 1 0 45540 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1636968456
transform 1 0 46644 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1
transform 1 0 47748 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1
transform 1 0 48300 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1636968456
transform 1 0 48484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1636968456
transform 1 0 49588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1636968456
transform 1 0 50692 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1636968456
transform 1 0 51796 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1
transform 1 0 52900 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1
transform 1 0 53452 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1636968456
transform 1 0 53636 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1636968456
transform 1 0 54740 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1636968456
transform 1 0 55844 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1636968456
transform 1 0 56948 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1
transform 1 0 58052 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1
transform 1 0 58604 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_617
timestamp 1636968456
transform 1 0 58788 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_629
timestamp 1636968456
transform 1 0 59892 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_641
timestamp 1636968456
transform 1 0 60996 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_653
timestamp 1636968456
transform 1 0 62100 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1
transform 1 0 63204 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1
transform 1 0 63756 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_673
timestamp 1636968456
transform 1 0 63940 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_685
timestamp 1636968456
transform 1 0 65044 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_697
timestamp 1636968456
transform 1 0 66148 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_709
timestamp 1636968456
transform 1 0 67252 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_721
timestamp 1
transform 1 0 68356 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_727
timestamp 1
transform 1 0 68908 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_729
timestamp 1636968456
transform 1 0 69092 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_741
timestamp 1636968456
transform 1 0 70196 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_753
timestamp 1636968456
transform 1 0 71300 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_765
timestamp 1636968456
transform 1 0 72404 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_777
timestamp 1
transform 1 0 73508 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_783
timestamp 1
transform 1 0 74060 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_785
timestamp 1636968456
transform 1 0 74244 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_797
timestamp 1636968456
transform 1 0 75348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_809
timestamp 1636968456
transform 1 0 76452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_821
timestamp 1
transform 1 0 77556 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1636968456
transform 1 0 2300 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1636968456
transform 1 0 3404 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1
transform 1 0 4508 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1636968456
transform 1 0 4692 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1636968456
transform 1 0 5796 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1636968456
transform 1 0 6900 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1636968456
transform 1 0 8004 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1
transform 1 0 9108 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1
transform 1 0 9660 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1636968456
transform 1 0 9844 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1636968456
transform 1 0 10948 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1636968456
transform 1 0 12052 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1636968456
transform 1 0 13156 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1
transform 1 0 14260 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1
transform 1 0 14812 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1636968456
transform 1 0 14996 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1636968456
transform 1 0 16100 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1636968456
transform 1 0 17204 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1636968456
transform 1 0 18308 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1
transform 1 0 19412 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1
transform 1 0 19964 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1636968456
transform 1 0 20148 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1636968456
transform 1 0 21252 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1636968456
transform 1 0 22356 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1636968456
transform 1 0 23460 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1
transform 1 0 24564 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1
transform 1 0 25116 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1636968456
transform 1 0 25300 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1636968456
transform 1 0 26404 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1636968456
transform 1 0 27508 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1636968456
transform 1 0 28612 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1
transform 1 0 29716 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1
transform 1 0 30268 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1636968456
transform 1 0 30452 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1636968456
transform 1 0 31556 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1636968456
transform 1 0 32660 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1636968456
transform 1 0 33764 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1
transform 1 0 34868 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1
transform 1 0 35420 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1636968456
transform 1 0 35604 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1636968456
transform 1 0 36708 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1636968456
transform 1 0 37812 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1636968456
transform 1 0 38916 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1
transform 1 0 40020 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1
transform 1 0 40572 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1636968456
transform 1 0 40756 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1636968456
transform 1 0 41860 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1636968456
transform 1 0 42964 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1636968456
transform 1 0 44068 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1
transform 1 0 45172 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1
transform 1 0 45724 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1636968456
transform 1 0 45908 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1636968456
transform 1 0 47012 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1636968456
transform 1 0 48116 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1636968456
transform 1 0 49220 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1
transform 1 0 50324 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1
transform 1 0 50876 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1636968456
transform 1 0 51060 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1636968456
transform 1 0 52164 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1636968456
transform 1 0 53268 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1636968456
transform 1 0 54372 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1
transform 1 0 55476 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1
transform 1 0 56028 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1636968456
transform 1 0 56212 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1636968456
transform 1 0 57316 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1636968456
transform 1 0 58420 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_625
timestamp 1636968456
transform 1 0 59524 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1
transform 1 0 60628 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1
transform 1 0 61180 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_645
timestamp 1636968456
transform 1 0 61364 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_657
timestamp 1636968456
transform 1 0 62468 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_669
timestamp 1636968456
transform 1 0 63572 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_681
timestamp 1636968456
transform 1 0 64676 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1
transform 1 0 65780 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1
transform 1 0 66332 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_701
timestamp 1636968456
transform 1 0 66516 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_713
timestamp 1636968456
transform 1 0 67620 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_725
timestamp 1636968456
transform 1 0 68724 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_737
timestamp 1636968456
transform 1 0 69828 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_749
timestamp 1
transform 1 0 70932 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_755
timestamp 1
transform 1 0 71484 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_757
timestamp 1636968456
transform 1 0 71668 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_769
timestamp 1636968456
transform 1 0 72772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_781
timestamp 1636968456
transform 1 0 73876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_793
timestamp 1636968456
transform 1 0 74980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_805
timestamp 1
transform 1 0 76084 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_811
timestamp 1
transform 1 0 76636 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_813
timestamp 1
transform 1 0 76820 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_821
timestamp 1
transform 1 0 77556 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1636968456
transform 1 0 2300 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1636968456
transform 1 0 3404 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1636968456
transform 1 0 4508 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1636968456
transform 1 0 5612 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1
transform 1 0 6716 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1636968456
transform 1 0 7268 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1636968456
transform 1 0 8372 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1636968456
transform 1 0 9476 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1636968456
transform 1 0 10580 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1
transform 1 0 11684 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1
transform 1 0 12236 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1636968456
transform 1 0 12420 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1636968456
transform 1 0 13524 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1636968456
transform 1 0 14628 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1636968456
transform 1 0 15732 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1
transform 1 0 16836 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1
transform 1 0 17388 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1636968456
transform 1 0 17572 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1636968456
transform 1 0 18676 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1636968456
transform 1 0 19780 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1636968456
transform 1 0 20884 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1
transform 1 0 21988 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1
transform 1 0 22540 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1636968456
transform 1 0 22724 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1636968456
transform 1 0 23828 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1636968456
transform 1 0 24932 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1636968456
transform 1 0 26036 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1
transform 1 0 27140 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1
transform 1 0 27692 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1636968456
transform 1 0 27876 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1636968456
transform 1 0 28980 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1636968456
transform 1 0 30084 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1636968456
transform 1 0 31188 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1
transform 1 0 32292 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1
transform 1 0 32844 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1636968456
transform 1 0 33028 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1636968456
transform 1 0 34132 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1636968456
transform 1 0 35236 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1636968456
transform 1 0 36340 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1
transform 1 0 37444 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1
transform 1 0 37996 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1636968456
transform 1 0 38180 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1636968456
transform 1 0 39284 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1636968456
transform 1 0 40388 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1636968456
transform 1 0 41492 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1
transform 1 0 42596 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1
transform 1 0 43148 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1636968456
transform 1 0 43332 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1636968456
transform 1 0 44436 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1636968456
transform 1 0 45540 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1636968456
transform 1 0 46644 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1
transform 1 0 47748 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1
transform 1 0 48300 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1636968456
transform 1 0 48484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1636968456
transform 1 0 49588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1636968456
transform 1 0 50692 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1636968456
transform 1 0 51796 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1
transform 1 0 52900 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1
transform 1 0 53452 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1636968456
transform 1 0 53636 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1636968456
transform 1 0 54740 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1636968456
transform 1 0 55844 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1636968456
transform 1 0 56948 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1
transform 1 0 58052 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1
transform 1 0 58604 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_617
timestamp 1636968456
transform 1 0 58788 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_629
timestamp 1636968456
transform 1 0 59892 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_641
timestamp 1636968456
transform 1 0 60996 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_653
timestamp 1636968456
transform 1 0 62100 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1
transform 1 0 63204 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1
transform 1 0 63756 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_673
timestamp 1636968456
transform 1 0 63940 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_685
timestamp 1636968456
transform 1 0 65044 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_697
timestamp 1636968456
transform 1 0 66148 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_709
timestamp 1636968456
transform 1 0 67252 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_721
timestamp 1
transform 1 0 68356 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_727
timestamp 1
transform 1 0 68908 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_729
timestamp 1636968456
transform 1 0 69092 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_741
timestamp 1636968456
transform 1 0 70196 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_753
timestamp 1636968456
transform 1 0 71300 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_765
timestamp 1636968456
transform 1 0 72404 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_777
timestamp 1
transform 1 0 73508 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_783
timestamp 1
transform 1 0 74060 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_785
timestamp 1636968456
transform 1 0 74244 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_797
timestamp 1636968456
transform 1 0 75348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_809
timestamp 1636968456
transform 1 0 76452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_95_821
timestamp 1
transform 1 0 77556 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1636968456
transform 1 0 2300 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1636968456
transform 1 0 3404 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1
transform 1 0 4508 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1636968456
transform 1 0 4692 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1636968456
transform 1 0 5796 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1636968456
transform 1 0 6900 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1636968456
transform 1 0 8004 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1
transform 1 0 9108 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1
transform 1 0 9660 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1636968456
transform 1 0 9844 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1636968456
transform 1 0 10948 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1636968456
transform 1 0 12052 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1636968456
transform 1 0 13156 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1
transform 1 0 14260 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1
transform 1 0 14812 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1636968456
transform 1 0 14996 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1636968456
transform 1 0 16100 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1636968456
transform 1 0 17204 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1636968456
transform 1 0 18308 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1
transform 1 0 19412 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1
transform 1 0 19964 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1636968456
transform 1 0 20148 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1636968456
transform 1 0 21252 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1636968456
transform 1 0 22356 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1636968456
transform 1 0 23460 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1
transform 1 0 24564 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1
transform 1 0 25116 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1636968456
transform 1 0 25300 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1636968456
transform 1 0 26404 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1636968456
transform 1 0 27508 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1636968456
transform 1 0 28612 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1
transform 1 0 29716 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1
transform 1 0 30268 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1636968456
transform 1 0 30452 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1636968456
transform 1 0 31556 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1636968456
transform 1 0 32660 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1636968456
transform 1 0 33764 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1
transform 1 0 34868 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1
transform 1 0 35420 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1636968456
transform 1 0 35604 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1636968456
transform 1 0 36708 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1636968456
transform 1 0 37812 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1636968456
transform 1 0 38916 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1
transform 1 0 40020 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1
transform 1 0 40572 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1636968456
transform 1 0 40756 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1636968456
transform 1 0 41860 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1636968456
transform 1 0 42964 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1636968456
transform 1 0 44068 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1
transform 1 0 45172 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1
transform 1 0 45724 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1636968456
transform 1 0 45908 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1636968456
transform 1 0 47012 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1636968456
transform 1 0 48116 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1636968456
transform 1 0 49220 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1
transform 1 0 50324 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1
transform 1 0 50876 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1636968456
transform 1 0 51060 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1636968456
transform 1 0 52164 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1636968456
transform 1 0 53268 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1636968456
transform 1 0 54372 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1
transform 1 0 55476 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1
transform 1 0 56028 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1636968456
transform 1 0 56212 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1636968456
transform 1 0 57316 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1636968456
transform 1 0 58420 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_625
timestamp 1636968456
transform 1 0 59524 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_637
timestamp 1
transform 1 0 60628 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_643
timestamp 1
transform 1 0 61180 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_645
timestamp 1636968456
transform 1 0 61364 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_657
timestamp 1636968456
transform 1 0 62468 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_669
timestamp 1636968456
transform 1 0 63572 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_681
timestamp 1636968456
transform 1 0 64676 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_693
timestamp 1
transform 1 0 65780 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_699
timestamp 1
transform 1 0 66332 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_701
timestamp 1636968456
transform 1 0 66516 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_713
timestamp 1636968456
transform 1 0 67620 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_725
timestamp 1636968456
transform 1 0 68724 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_737
timestamp 1636968456
transform 1 0 69828 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_749
timestamp 1
transform 1 0 70932 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_755
timestamp 1
transform 1 0 71484 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_757
timestamp 1636968456
transform 1 0 71668 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_769
timestamp 1636968456
transform 1 0 72772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_781
timestamp 1636968456
transform 1 0 73876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_793
timestamp 1636968456
transform 1 0 74980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_805
timestamp 1
transform 1 0 76084 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_811
timestamp 1
transform 1 0 76636 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_813
timestamp 1
transform 1 0 76820 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_821
timestamp 1
transform 1 0 77556 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1636968456
transform 1 0 2300 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1636968456
transform 1 0 3404 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1636968456
transform 1 0 4508 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1636968456
transform 1 0 5612 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1
transform 1 0 6716 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1
transform 1 0 7084 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1636968456
transform 1 0 7268 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1636968456
transform 1 0 8372 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1636968456
transform 1 0 9476 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1636968456
transform 1 0 10580 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1
transform 1 0 11684 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1
transform 1 0 12236 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1636968456
transform 1 0 12420 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1636968456
transform 1 0 13524 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1636968456
transform 1 0 14628 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1636968456
transform 1 0 15732 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1
transform 1 0 16836 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1
transform 1 0 17388 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1636968456
transform 1 0 17572 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1636968456
transform 1 0 18676 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1636968456
transform 1 0 19780 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1636968456
transform 1 0 20884 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1
transform 1 0 21988 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1
transform 1 0 22540 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1636968456
transform 1 0 22724 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1636968456
transform 1 0 23828 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1636968456
transform 1 0 24932 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1636968456
transform 1 0 26036 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1
transform 1 0 27140 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1
transform 1 0 27692 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1636968456
transform 1 0 27876 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1636968456
transform 1 0 28980 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1636968456
transform 1 0 30084 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1636968456
transform 1 0 31188 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1
transform 1 0 32292 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1
transform 1 0 32844 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1636968456
transform 1 0 33028 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1636968456
transform 1 0 34132 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1636968456
transform 1 0 35236 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1636968456
transform 1 0 36340 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1
transform 1 0 37444 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1
transform 1 0 37996 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1636968456
transform 1 0 38180 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1636968456
transform 1 0 39284 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1636968456
transform 1 0 40388 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1636968456
transform 1 0 41492 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1
transform 1 0 42596 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1
transform 1 0 43148 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1636968456
transform 1 0 43332 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1636968456
transform 1 0 44436 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1636968456
transform 1 0 45540 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1636968456
transform 1 0 46644 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1
transform 1 0 47748 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1
transform 1 0 48300 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1636968456
transform 1 0 48484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1636968456
transform 1 0 49588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1636968456
transform 1 0 50692 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1636968456
transform 1 0 51796 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1
transform 1 0 52900 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1
transform 1 0 53452 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1636968456
transform 1 0 53636 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1636968456
transform 1 0 54740 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1636968456
transform 1 0 55844 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1636968456
transform 1 0 56948 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1
transform 1 0 58052 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1
transform 1 0 58604 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_617
timestamp 1636968456
transform 1 0 58788 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_629
timestamp 1636968456
transform 1 0 59892 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_641
timestamp 1636968456
transform 1 0 60996 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_653
timestamp 1636968456
transform 1 0 62100 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_665
timestamp 1
transform 1 0 63204 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_671
timestamp 1
transform 1 0 63756 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_673
timestamp 1636968456
transform 1 0 63940 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_685
timestamp 1636968456
transform 1 0 65044 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_697
timestamp 1636968456
transform 1 0 66148 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_709
timestamp 1636968456
transform 1 0 67252 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_721
timestamp 1
transform 1 0 68356 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_727
timestamp 1
transform 1 0 68908 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_729
timestamp 1636968456
transform 1 0 69092 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_741
timestamp 1636968456
transform 1 0 70196 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_753
timestamp 1636968456
transform 1 0 71300 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_765
timestamp 1636968456
transform 1 0 72404 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_777
timestamp 1
transform 1 0 73508 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_783
timestamp 1
transform 1 0 74060 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_785
timestamp 1636968456
transform 1 0 74244 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_797
timestamp 1636968456
transform 1 0 75348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_809
timestamp 1636968456
transform 1 0 76452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_821
timestamp 1
transform 1 0 77556 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1636968456
transform 1 0 2300 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1636968456
transform 1 0 3404 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1
transform 1 0 4508 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1636968456
transform 1 0 4692 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1636968456
transform 1 0 5796 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1636968456
transform 1 0 6900 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1636968456
transform 1 0 8004 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1
transform 1 0 9108 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1
transform 1 0 9660 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1636968456
transform 1 0 9844 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1636968456
transform 1 0 10948 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1636968456
transform 1 0 12052 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1636968456
transform 1 0 13156 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1
transform 1 0 14260 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1
transform 1 0 14812 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1636968456
transform 1 0 14996 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1636968456
transform 1 0 16100 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1636968456
transform 1 0 17204 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1636968456
transform 1 0 18308 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1
transform 1 0 19412 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1
transform 1 0 19964 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1636968456
transform 1 0 20148 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1636968456
transform 1 0 21252 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1636968456
transform 1 0 22356 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1636968456
transform 1 0 23460 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1
transform 1 0 24564 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1
transform 1 0 25116 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1636968456
transform 1 0 25300 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1636968456
transform 1 0 26404 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1636968456
transform 1 0 27508 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1636968456
transform 1 0 28612 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1
transform 1 0 29716 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1
transform 1 0 30268 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1636968456
transform 1 0 30452 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1636968456
transform 1 0 31556 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1636968456
transform 1 0 32660 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1636968456
transform 1 0 33764 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1
transform 1 0 34868 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1
transform 1 0 35420 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1636968456
transform 1 0 35604 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1636968456
transform 1 0 36708 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1636968456
transform 1 0 37812 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1636968456
transform 1 0 38916 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1
transform 1 0 40020 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1
transform 1 0 40572 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1636968456
transform 1 0 40756 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1636968456
transform 1 0 41860 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1636968456
transform 1 0 42964 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1636968456
transform 1 0 44068 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1
transform 1 0 45172 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1
transform 1 0 45724 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1636968456
transform 1 0 45908 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1636968456
transform 1 0 47012 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1636968456
transform 1 0 48116 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1636968456
transform 1 0 49220 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1
transform 1 0 50324 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1
transform 1 0 50876 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1636968456
transform 1 0 51060 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1636968456
transform 1 0 52164 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1636968456
transform 1 0 53268 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1636968456
transform 1 0 54372 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1
transform 1 0 55476 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1
transform 1 0 56028 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1636968456
transform 1 0 56212 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1636968456
transform 1 0 57316 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1636968456
transform 1 0 58420 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_625
timestamp 1636968456
transform 1 0 59524 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_637
timestamp 1
transform 1 0 60628 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_643
timestamp 1
transform 1 0 61180 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_645
timestamp 1636968456
transform 1 0 61364 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_657
timestamp 1636968456
transform 1 0 62468 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_669
timestamp 1636968456
transform 1 0 63572 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_681
timestamp 1636968456
transform 1 0 64676 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_693
timestamp 1
transform 1 0 65780 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_699
timestamp 1
transform 1 0 66332 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_701
timestamp 1636968456
transform 1 0 66516 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_713
timestamp 1636968456
transform 1 0 67620 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_725
timestamp 1636968456
transform 1 0 68724 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_737
timestamp 1636968456
transform 1 0 69828 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_749
timestamp 1
transform 1 0 70932 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_755
timestamp 1
transform 1 0 71484 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_757
timestamp 1636968456
transform 1 0 71668 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_769
timestamp 1636968456
transform 1 0 72772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_781
timestamp 1636968456
transform 1 0 73876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_793
timestamp 1636968456
transform 1 0 74980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_805
timestamp 1
transform 1 0 76084 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_811
timestamp 1
transform 1 0 76636 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_813
timestamp 1
transform 1 0 76820 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_821
timestamp 1
transform 1 0 77556 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1636968456
transform 1 0 2300 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1636968456
transform 1 0 3404 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1636968456
transform 1 0 4508 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1636968456
transform 1 0 5612 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1
transform 1 0 6716 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1
transform 1 0 7084 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1636968456
transform 1 0 7268 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1636968456
transform 1 0 8372 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1636968456
transform 1 0 9476 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1636968456
transform 1 0 10580 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1
transform 1 0 11684 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1
transform 1 0 12236 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1636968456
transform 1 0 12420 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1636968456
transform 1 0 13524 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1636968456
transform 1 0 14628 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1636968456
transform 1 0 15732 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1
transform 1 0 16836 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1
transform 1 0 17388 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1636968456
transform 1 0 17572 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1636968456
transform 1 0 18676 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1636968456
transform 1 0 19780 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1636968456
transform 1 0 20884 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1
transform 1 0 21988 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1
transform 1 0 22540 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1636968456
transform 1 0 22724 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1636968456
transform 1 0 23828 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1636968456
transform 1 0 24932 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1636968456
transform 1 0 26036 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1
transform 1 0 27140 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1
transform 1 0 27692 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1636968456
transform 1 0 27876 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1636968456
transform 1 0 28980 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1636968456
transform 1 0 30084 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1636968456
transform 1 0 31188 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1
transform 1 0 32292 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1
transform 1 0 32844 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1636968456
transform 1 0 33028 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1636968456
transform 1 0 34132 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1636968456
transform 1 0 35236 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1636968456
transform 1 0 36340 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1
transform 1 0 37444 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1
transform 1 0 37996 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1636968456
transform 1 0 38180 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1636968456
transform 1 0 39284 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1636968456
transform 1 0 40388 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1636968456
transform 1 0 41492 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1
transform 1 0 42596 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1
transform 1 0 43148 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1636968456
transform 1 0 43332 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1636968456
transform 1 0 44436 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1636968456
transform 1 0 45540 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1636968456
transform 1 0 46644 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1
transform 1 0 47748 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1
transform 1 0 48300 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1636968456
transform 1 0 48484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1636968456
transform 1 0 49588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1636968456
transform 1 0 50692 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1636968456
transform 1 0 51796 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1
transform 1 0 52900 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1
transform 1 0 53452 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1636968456
transform 1 0 53636 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1636968456
transform 1 0 54740 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1636968456
transform 1 0 55844 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1636968456
transform 1 0 56948 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1
transform 1 0 58052 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1
transform 1 0 58604 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_617
timestamp 1636968456
transform 1 0 58788 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_629
timestamp 1636968456
transform 1 0 59892 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_641
timestamp 1636968456
transform 1 0 60996 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_653
timestamp 1636968456
transform 1 0 62100 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_665
timestamp 1
transform 1 0 63204 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1
transform 1 0 63756 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_673
timestamp 1636968456
transform 1 0 63940 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_685
timestamp 1636968456
transform 1 0 65044 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_697
timestamp 1636968456
transform 1 0 66148 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_709
timestamp 1636968456
transform 1 0 67252 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_721
timestamp 1
transform 1 0 68356 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_727
timestamp 1
transform 1 0 68908 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_729
timestamp 1636968456
transform 1 0 69092 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_741
timestamp 1636968456
transform 1 0 70196 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_753
timestamp 1636968456
transform 1 0 71300 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_765
timestamp 1636968456
transform 1 0 72404 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_777
timestamp 1
transform 1 0 73508 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_783
timestamp 1
transform 1 0 74060 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_785
timestamp 1636968456
transform 1 0 74244 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_797
timestamp 1636968456
transform 1 0 75348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_809
timestamp 1636968456
transform 1 0 76452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_821
timestamp 1
transform 1 0 77556 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1636968456
transform 1 0 2300 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1636968456
transform 1 0 3404 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1
transform 1 0 4508 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1636968456
transform 1 0 4692 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1636968456
transform 1 0 5796 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1636968456
transform 1 0 6900 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1636968456
transform 1 0 8004 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1
transform 1 0 9108 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1
transform 1 0 9660 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1636968456
transform 1 0 9844 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1636968456
transform 1 0 10948 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1636968456
transform 1 0 12052 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1636968456
transform 1 0 13156 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1
transform 1 0 14260 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1
transform 1 0 14812 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1636968456
transform 1 0 14996 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1636968456
transform 1 0 16100 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1636968456
transform 1 0 17204 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1636968456
transform 1 0 18308 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1
transform 1 0 19412 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1
transform 1 0 19964 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1636968456
transform 1 0 20148 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1636968456
transform 1 0 21252 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1636968456
transform 1 0 22356 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1636968456
transform 1 0 23460 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1
transform 1 0 24564 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1
transform 1 0 25116 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1636968456
transform 1 0 25300 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1636968456
transform 1 0 26404 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1636968456
transform 1 0 27508 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1636968456
transform 1 0 28612 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1
transform 1 0 29716 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1
transform 1 0 30268 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1636968456
transform 1 0 30452 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1636968456
transform 1 0 31556 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1636968456
transform 1 0 32660 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1636968456
transform 1 0 33764 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1
transform 1 0 34868 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1
transform 1 0 35420 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1636968456
transform 1 0 35604 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1636968456
transform 1 0 36708 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1636968456
transform 1 0 37812 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1636968456
transform 1 0 38916 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1
transform 1 0 40020 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1
transform 1 0 40572 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1636968456
transform 1 0 40756 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1636968456
transform 1 0 41860 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1636968456
transform 1 0 42964 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1636968456
transform 1 0 44068 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1
transform 1 0 45172 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1
transform 1 0 45724 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1636968456
transform 1 0 45908 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1636968456
transform 1 0 47012 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1636968456
transform 1 0 48116 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1636968456
transform 1 0 49220 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1
transform 1 0 50324 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1
transform 1 0 50876 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1636968456
transform 1 0 51060 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1636968456
transform 1 0 52164 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1636968456
transform 1 0 53268 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1636968456
transform 1 0 54372 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1
transform 1 0 55476 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1
transform 1 0 56028 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1636968456
transform 1 0 56212 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1636968456
transform 1 0 57316 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1636968456
transform 1 0 58420 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_625
timestamp 1636968456
transform 1 0 59524 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_637
timestamp 1
transform 1 0 60628 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_643
timestamp 1
transform 1 0 61180 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_645
timestamp 1636968456
transform 1 0 61364 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_657
timestamp 1636968456
transform 1 0 62468 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_669
timestamp 1636968456
transform 1 0 63572 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_681
timestamp 1636968456
transform 1 0 64676 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_693
timestamp 1
transform 1 0 65780 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_699
timestamp 1
transform 1 0 66332 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_701
timestamp 1636968456
transform 1 0 66516 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_713
timestamp 1636968456
transform 1 0 67620 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_725
timestamp 1636968456
transform 1 0 68724 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_737
timestamp 1636968456
transform 1 0 69828 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_749
timestamp 1
transform 1 0 70932 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_755
timestamp 1
transform 1 0 71484 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_757
timestamp 1636968456
transform 1 0 71668 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_769
timestamp 1636968456
transform 1 0 72772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_781
timestamp 1636968456
transform 1 0 73876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_793
timestamp 1636968456
transform 1 0 74980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_805
timestamp 1
transform 1 0 76084 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_811
timestamp 1
transform 1 0 76636 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_813
timestamp 1
transform 1 0 76820 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_821
timestamp 1
transform 1 0 77556 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1636968456
transform 1 0 2300 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1636968456
transform 1 0 3404 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_27
timestamp 1636968456
transform 1 0 4508 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_39
timestamp 1636968456
transform 1 0 5612 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1
transform 1 0 6716 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1
transform 1 0 7084 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1636968456
transform 1 0 7268 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1636968456
transform 1 0 8372 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_81
timestamp 1636968456
transform 1 0 9476 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_93
timestamp 1636968456
transform 1 0 10580 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1
transform 1 0 11684 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1
transform 1 0 12236 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1636968456
transform 1 0 12420 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1636968456
transform 1 0 13524 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_137
timestamp 1636968456
transform 1 0 14628 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_149
timestamp 1636968456
transform 1 0 15732 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_161
timestamp 1
transform 1 0 16836 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1
transform 1 0 17388 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1636968456
transform 1 0 17572 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1636968456
transform 1 0 18676 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_193
timestamp 1636968456
transform 1 0 19780 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_205
timestamp 1636968456
transform 1 0 20884 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_217
timestamp 1
transform 1 0 21988 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1
transform 1 0 22540 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1636968456
transform 1 0 22724 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1636968456
transform 1 0 23828 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_249
timestamp 1636968456
transform 1 0 24932 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_261
timestamp 1636968456
transform 1 0 26036 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1
transform 1 0 27140 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1
transform 1 0 27692 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1636968456
transform 1 0 27876 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1636968456
transform 1 0 28980 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_305
timestamp 1636968456
transform 1 0 30084 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_317
timestamp 1636968456
transform 1 0 31188 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_329
timestamp 1
transform 1 0 32292 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_335
timestamp 1
transform 1 0 32844 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1636968456
transform 1 0 33028 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1636968456
transform 1 0 34132 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_361
timestamp 1636968456
transform 1 0 35236 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_373
timestamp 1636968456
transform 1 0 36340 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_385
timestamp 1
transform 1 0 37444 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_391
timestamp 1
transform 1 0 37996 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1636968456
transform 1 0 38180 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1636968456
transform 1 0 39284 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_417
timestamp 1636968456
transform 1 0 40388 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_429
timestamp 1636968456
transform 1 0 41492 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1
transform 1 0 42596 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1
transform 1 0 43148 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1636968456
transform 1 0 43332 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1636968456
transform 1 0 44436 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_473
timestamp 1636968456
transform 1 0 45540 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_485
timestamp 1636968456
transform 1 0 46644 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1
transform 1 0 47748 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1
transform 1 0 48300 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1636968456
transform 1 0 48484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1636968456
transform 1 0 49588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_529
timestamp 1636968456
transform 1 0 50692 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_541
timestamp 1636968456
transform 1 0 51796 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_553
timestamp 1
transform 1 0 52900 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1
transform 1 0 53452 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1636968456
transform 1 0 53636 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1636968456
transform 1 0 54740 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_585
timestamp 1636968456
transform 1 0 55844 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_597
timestamp 1636968456
transform 1 0 56948 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_609
timestamp 1
transform 1 0 58052 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1
transform 1 0 58604 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_617
timestamp 1636968456
transform 1 0 58788 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_629
timestamp 1636968456
transform 1 0 59892 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_641
timestamp 1636968456
transform 1 0 60996 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_653
timestamp 1636968456
transform 1 0 62100 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_665
timestamp 1
transform 1 0 63204 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_671
timestamp 1
transform 1 0 63756 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_673
timestamp 1636968456
transform 1 0 63940 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_685
timestamp 1636968456
transform 1 0 65044 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_697
timestamp 1636968456
transform 1 0 66148 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_709
timestamp 1636968456
transform 1 0 67252 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_721
timestamp 1
transform 1 0 68356 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_727
timestamp 1
transform 1 0 68908 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_729
timestamp 1636968456
transform 1 0 69092 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_741
timestamp 1636968456
transform 1 0 70196 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_753
timestamp 1636968456
transform 1 0 71300 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_765
timestamp 1636968456
transform 1 0 72404 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_777
timestamp 1
transform 1 0 73508 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_783
timestamp 1
transform 1 0 74060 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_785
timestamp 1636968456
transform 1 0 74244 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_797
timestamp 1636968456
transform 1 0 75348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_809
timestamp 1636968456
transform 1 0 76452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_821
timestamp 1
transform 1 0 77556 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_3
timestamp 1636968456
transform 1 0 2300 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_15
timestamp 1636968456
transform 1 0 3404 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1
transform 1 0 4508 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1636968456
transform 1 0 4692 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1636968456
transform 1 0 5796 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1636968456
transform 1 0 6900 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_65
timestamp 1636968456
transform 1 0 8004 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1
transform 1 0 9108 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1
transform 1 0 9660 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_85
timestamp 1636968456
transform 1 0 9844 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_97
timestamp 1636968456
transform 1 0 10948 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_109
timestamp 1636968456
transform 1 0 12052 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_121
timestamp 1636968456
transform 1 0 13156 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1
transform 1 0 14260 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1
transform 1 0 14812 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_141
timestamp 1636968456
transform 1 0 14996 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_153
timestamp 1636968456
transform 1 0 16100 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_165
timestamp 1636968456
transform 1 0 17204 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_177
timestamp 1636968456
transform 1 0 18308 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_189
timestamp 1
transform 1 0 19412 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1
transform 1 0 19964 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_197
timestamp 1636968456
transform 1 0 20148 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_209
timestamp 1636968456
transform 1 0 21252 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_221
timestamp 1636968456
transform 1 0 22356 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_233
timestamp 1636968456
transform 1 0 23460 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_245
timestamp 1
transform 1 0 24564 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_251
timestamp 1
transform 1 0 25116 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_253
timestamp 1636968456
transform 1 0 25300 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_265
timestamp 1636968456
transform 1 0 26404 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_277
timestamp 1636968456
transform 1 0 27508 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_289
timestamp 1636968456
transform 1 0 28612 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_301
timestamp 1
transform 1 0 29716 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_307
timestamp 1
transform 1 0 30268 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_309
timestamp 1636968456
transform 1 0 30452 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_321
timestamp 1636968456
transform 1 0 31556 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_333
timestamp 1636968456
transform 1 0 32660 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_345
timestamp 1636968456
transform 1 0 33764 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_357
timestamp 1
transform 1 0 34868 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_363
timestamp 1
transform 1 0 35420 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_365
timestamp 1636968456
transform 1 0 35604 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_377
timestamp 1636968456
transform 1 0 36708 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_389
timestamp 1636968456
transform 1 0 37812 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_401
timestamp 1636968456
transform 1 0 38916 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_413
timestamp 1
transform 1 0 40020 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_419
timestamp 1
transform 1 0 40572 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_421
timestamp 1636968456
transform 1 0 40756 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_433
timestamp 1636968456
transform 1 0 41860 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_445
timestamp 1636968456
transform 1 0 42964 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_457
timestamp 1636968456
transform 1 0 44068 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_469
timestamp 1
transform 1 0 45172 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_475
timestamp 1
transform 1 0 45724 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_477
timestamp 1636968456
transform 1 0 45908 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_489
timestamp 1636968456
transform 1 0 47012 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_501
timestamp 1636968456
transform 1 0 48116 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_513
timestamp 1636968456
transform 1 0 49220 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_525
timestamp 1
transform 1 0 50324 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_531
timestamp 1
transform 1 0 50876 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_533
timestamp 1636968456
transform 1 0 51060 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_545
timestamp 1636968456
transform 1 0 52164 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_557
timestamp 1636968456
transform 1 0 53268 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_569
timestamp 1636968456
transform 1 0 54372 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_581
timestamp 1
transform 1 0 55476 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_587
timestamp 1
transform 1 0 56028 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_589
timestamp 1636968456
transform 1 0 56212 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_601
timestamp 1636968456
transform 1 0 57316 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_613
timestamp 1636968456
transform 1 0 58420 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_625
timestamp 1636968456
transform 1 0 59524 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_637
timestamp 1
transform 1 0 60628 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_643
timestamp 1
transform 1 0 61180 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_645
timestamp 1636968456
transform 1 0 61364 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_657
timestamp 1636968456
transform 1 0 62468 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_669
timestamp 1636968456
transform 1 0 63572 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_681
timestamp 1636968456
transform 1 0 64676 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_693
timestamp 1
transform 1 0 65780 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_699
timestamp 1
transform 1 0 66332 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_701
timestamp 1636968456
transform 1 0 66516 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_713
timestamp 1636968456
transform 1 0 67620 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_725
timestamp 1636968456
transform 1 0 68724 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_737
timestamp 1636968456
transform 1 0 69828 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_749
timestamp 1
transform 1 0 70932 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_755
timestamp 1
transform 1 0 71484 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_757
timestamp 1636968456
transform 1 0 71668 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_769
timestamp 1636968456
transform 1 0 72772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_781
timestamp 1636968456
transform 1 0 73876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_793
timestamp 1636968456
transform 1 0 74980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_805
timestamp 1
transform 1 0 76084 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_811
timestamp 1
transform 1 0 76636 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_813
timestamp 1
transform 1 0 76820 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_102_821
timestamp 1
transform 1 0 77556 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_3
timestamp 1636968456
transform 1 0 2300 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_15
timestamp 1636968456
transform 1 0 3404 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_27
timestamp 1636968456
transform 1 0 4508 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_39
timestamp 1636968456
transform 1 0 5612 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_51
timestamp 1
transform 1 0 6716 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1
transform 1 0 7084 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1636968456
transform 1 0 7268 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_69
timestamp 1636968456
transform 1 0 8372 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_81
timestamp 1636968456
transform 1 0 9476 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_93
timestamp 1636968456
transform 1 0 10580 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1
transform 1 0 11684 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1
transform 1 0 12236 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_113
timestamp 1636968456
transform 1 0 12420 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_125
timestamp 1636968456
transform 1 0 13524 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_137
timestamp 1636968456
transform 1 0 14628 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_149
timestamp 1636968456
transform 1 0 15732 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_161
timestamp 1
transform 1 0 16836 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_167
timestamp 1
transform 1 0 17388 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_169
timestamp 1636968456
transform 1 0 17572 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_181
timestamp 1636968456
transform 1 0 18676 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_193
timestamp 1636968456
transform 1 0 19780 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_205
timestamp 1636968456
transform 1 0 20884 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_217
timestamp 1
transform 1 0 21988 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_223
timestamp 1
transform 1 0 22540 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_225
timestamp 1636968456
transform 1 0 22724 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_237
timestamp 1636968456
transform 1 0 23828 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_249
timestamp 1636968456
transform 1 0 24932 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_261
timestamp 1636968456
transform 1 0 26036 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_273
timestamp 1
transform 1 0 27140 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_279
timestamp 1
transform 1 0 27692 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_281
timestamp 1636968456
transform 1 0 27876 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_293
timestamp 1636968456
transform 1 0 28980 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_305
timestamp 1636968456
transform 1 0 30084 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_317
timestamp 1636968456
transform 1 0 31188 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_329
timestamp 1
transform 1 0 32292 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_335
timestamp 1
transform 1 0 32844 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_337
timestamp 1636968456
transform 1 0 33028 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_349
timestamp 1636968456
transform 1 0 34132 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_361
timestamp 1636968456
transform 1 0 35236 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_373
timestamp 1636968456
transform 1 0 36340 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_385
timestamp 1
transform 1 0 37444 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_391
timestamp 1
transform 1 0 37996 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_393
timestamp 1636968456
transform 1 0 38180 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_405
timestamp 1636968456
transform 1 0 39284 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_417
timestamp 1636968456
transform 1 0 40388 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_429
timestamp 1636968456
transform 1 0 41492 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_441
timestamp 1
transform 1 0 42596 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_447
timestamp 1
transform 1 0 43148 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_449
timestamp 1636968456
transform 1 0 43332 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_461
timestamp 1636968456
transform 1 0 44436 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_473
timestamp 1636968456
transform 1 0 45540 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_485
timestamp 1636968456
transform 1 0 46644 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_497
timestamp 1
transform 1 0 47748 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_503
timestamp 1
transform 1 0 48300 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_505
timestamp 1636968456
transform 1 0 48484 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_517
timestamp 1636968456
transform 1 0 49588 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_529
timestamp 1636968456
transform 1 0 50692 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_541
timestamp 1636968456
transform 1 0 51796 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_553
timestamp 1
transform 1 0 52900 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_559
timestamp 1
transform 1 0 53452 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_561
timestamp 1636968456
transform 1 0 53636 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_573
timestamp 1636968456
transform 1 0 54740 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_585
timestamp 1636968456
transform 1 0 55844 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_597
timestamp 1636968456
transform 1 0 56948 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_609
timestamp 1
transform 1 0 58052 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_615
timestamp 1
transform 1 0 58604 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_617
timestamp 1636968456
transform 1 0 58788 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_629
timestamp 1636968456
transform 1 0 59892 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_641
timestamp 1636968456
transform 1 0 60996 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_653
timestamp 1636968456
transform 1 0 62100 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_665
timestamp 1
transform 1 0 63204 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_671
timestamp 1
transform 1 0 63756 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_673
timestamp 1636968456
transform 1 0 63940 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_685
timestamp 1636968456
transform 1 0 65044 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_697
timestamp 1636968456
transform 1 0 66148 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_709
timestamp 1636968456
transform 1 0 67252 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_721
timestamp 1
transform 1 0 68356 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_727
timestamp 1
transform 1 0 68908 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_729
timestamp 1636968456
transform 1 0 69092 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_741
timestamp 1636968456
transform 1 0 70196 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_753
timestamp 1636968456
transform 1 0 71300 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_765
timestamp 1636968456
transform 1 0 72404 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_777
timestamp 1
transform 1 0 73508 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_783
timestamp 1
transform 1 0 74060 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_785
timestamp 1636968456
transform 1 0 74244 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_797
timestamp 1636968456
transform 1 0 75348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_809
timestamp 1636968456
transform 1 0 76452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_103_821
timestamp 1
transform 1 0 77556 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_3
timestamp 1636968456
transform 1 0 2300 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_15
timestamp 1636968456
transform 1 0 3404 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1
transform 1 0 4508 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1636968456
transform 1 0 4692 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1636968456
transform 1 0 5796 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1636968456
transform 1 0 6900 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_65
timestamp 1636968456
transform 1 0 8004 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1
transform 1 0 9108 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1
transform 1 0 9660 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_85
timestamp 1636968456
transform 1 0 9844 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_97
timestamp 1636968456
transform 1 0 10948 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_109
timestamp 1636968456
transform 1 0 12052 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_121
timestamp 1636968456
transform 1 0 13156 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1
transform 1 0 14260 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1
transform 1 0 14812 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_141
timestamp 1636968456
transform 1 0 14996 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_153
timestamp 1636968456
transform 1 0 16100 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_165
timestamp 1636968456
transform 1 0 17204 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_177
timestamp 1636968456
transform 1 0 18308 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_189
timestamp 1
transform 1 0 19412 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_195
timestamp 1
transform 1 0 19964 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_197
timestamp 1636968456
transform 1 0 20148 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_209
timestamp 1636968456
transform 1 0 21252 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_221
timestamp 1636968456
transform 1 0 22356 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_233
timestamp 1636968456
transform 1 0 23460 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_245
timestamp 1
transform 1 0 24564 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_251
timestamp 1
transform 1 0 25116 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_253
timestamp 1636968456
transform 1 0 25300 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_265
timestamp 1636968456
transform 1 0 26404 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_277
timestamp 1636968456
transform 1 0 27508 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_289
timestamp 1636968456
transform 1 0 28612 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_301
timestamp 1
transform 1 0 29716 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_307
timestamp 1
transform 1 0 30268 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_309
timestamp 1636968456
transform 1 0 30452 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_321
timestamp 1636968456
transform 1 0 31556 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_333
timestamp 1636968456
transform 1 0 32660 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_345
timestamp 1636968456
transform 1 0 33764 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_357
timestamp 1
transform 1 0 34868 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_363
timestamp 1
transform 1 0 35420 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_365
timestamp 1636968456
transform 1 0 35604 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_377
timestamp 1636968456
transform 1 0 36708 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_389
timestamp 1636968456
transform 1 0 37812 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_401
timestamp 1636968456
transform 1 0 38916 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_413
timestamp 1
transform 1 0 40020 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_419
timestamp 1
transform 1 0 40572 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_421
timestamp 1636968456
transform 1 0 40756 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_433
timestamp 1636968456
transform 1 0 41860 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_445
timestamp 1636968456
transform 1 0 42964 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_457
timestamp 1636968456
transform 1 0 44068 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_469
timestamp 1
transform 1 0 45172 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_475
timestamp 1
transform 1 0 45724 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_477
timestamp 1636968456
transform 1 0 45908 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_489
timestamp 1636968456
transform 1 0 47012 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_501
timestamp 1636968456
transform 1 0 48116 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_513
timestamp 1636968456
transform 1 0 49220 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_525
timestamp 1
transform 1 0 50324 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_531
timestamp 1
transform 1 0 50876 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_533
timestamp 1636968456
transform 1 0 51060 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_545
timestamp 1636968456
transform 1 0 52164 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_557
timestamp 1636968456
transform 1 0 53268 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_569
timestamp 1636968456
transform 1 0 54372 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_581
timestamp 1
transform 1 0 55476 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_587
timestamp 1
transform 1 0 56028 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_589
timestamp 1636968456
transform 1 0 56212 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_601
timestamp 1636968456
transform 1 0 57316 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_613
timestamp 1636968456
transform 1 0 58420 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_625
timestamp 1636968456
transform 1 0 59524 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_637
timestamp 1
transform 1 0 60628 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_643
timestamp 1
transform 1 0 61180 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_645
timestamp 1636968456
transform 1 0 61364 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_657
timestamp 1636968456
transform 1 0 62468 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_669
timestamp 1636968456
transform 1 0 63572 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_681
timestamp 1636968456
transform 1 0 64676 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_693
timestamp 1
transform 1 0 65780 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_699
timestamp 1
transform 1 0 66332 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_701
timestamp 1636968456
transform 1 0 66516 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_713
timestamp 1636968456
transform 1 0 67620 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_725
timestamp 1636968456
transform 1 0 68724 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_737
timestamp 1636968456
transform 1 0 69828 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_749
timestamp 1
transform 1 0 70932 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_755
timestamp 1
transform 1 0 71484 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_757
timestamp 1636968456
transform 1 0 71668 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_769
timestamp 1636968456
transform 1 0 72772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_781
timestamp 1636968456
transform 1 0 73876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_793
timestamp 1636968456
transform 1 0 74980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_805
timestamp 1
transform 1 0 76084 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_811
timestamp 1
transform 1 0 76636 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_813
timestamp 1
transform 1 0 76820 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_821
timestamp 1
transform 1 0 77556 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_3
timestamp 1636968456
transform 1 0 2300 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_15
timestamp 1636968456
transform 1 0 3404 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_27
timestamp 1636968456
transform 1 0 4508 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_39
timestamp 1636968456
transform 1 0 5612 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1
transform 1 0 6716 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1
transform 1 0 7084 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1636968456
transform 1 0 7268 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_69
timestamp 1636968456
transform 1 0 8372 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_81
timestamp 1636968456
transform 1 0 9476 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_93
timestamp 1636968456
transform 1 0 10580 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1
transform 1 0 11684 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1
transform 1 0 12236 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_113
timestamp 1636968456
transform 1 0 12420 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_125
timestamp 1636968456
transform 1 0 13524 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_137
timestamp 1636968456
transform 1 0 14628 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_149
timestamp 1636968456
transform 1 0 15732 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1
transform 1 0 16836 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1
transform 1 0 17388 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_169
timestamp 1636968456
transform 1 0 17572 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_181
timestamp 1636968456
transform 1 0 18676 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_193
timestamp 1636968456
transform 1 0 19780 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_205
timestamp 1636968456
transform 1 0 20884 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_217
timestamp 1
transform 1 0 21988 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_223
timestamp 1
transform 1 0 22540 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_225
timestamp 1636968456
transform 1 0 22724 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_237
timestamp 1636968456
transform 1 0 23828 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_249
timestamp 1636968456
transform 1 0 24932 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_261
timestamp 1636968456
transform 1 0 26036 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_273
timestamp 1
transform 1 0 27140 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_279
timestamp 1
transform 1 0 27692 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_281
timestamp 1636968456
transform 1 0 27876 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_293
timestamp 1636968456
transform 1 0 28980 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_305
timestamp 1636968456
transform 1 0 30084 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_317
timestamp 1636968456
transform 1 0 31188 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_329
timestamp 1
transform 1 0 32292 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_335
timestamp 1
transform 1 0 32844 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_337
timestamp 1636968456
transform 1 0 33028 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_349
timestamp 1636968456
transform 1 0 34132 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_361
timestamp 1636968456
transform 1 0 35236 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_373
timestamp 1636968456
transform 1 0 36340 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_385
timestamp 1
transform 1 0 37444 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_391
timestamp 1
transform 1 0 37996 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_393
timestamp 1636968456
transform 1 0 38180 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_405
timestamp 1636968456
transform 1 0 39284 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_417
timestamp 1636968456
transform 1 0 40388 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_429
timestamp 1636968456
transform 1 0 41492 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_441
timestamp 1
transform 1 0 42596 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_447
timestamp 1
transform 1 0 43148 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_449
timestamp 1636968456
transform 1 0 43332 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_461
timestamp 1636968456
transform 1 0 44436 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_473
timestamp 1636968456
transform 1 0 45540 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_485
timestamp 1636968456
transform 1 0 46644 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_497
timestamp 1
transform 1 0 47748 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_503
timestamp 1
transform 1 0 48300 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_505
timestamp 1636968456
transform 1 0 48484 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_517
timestamp 1636968456
transform 1 0 49588 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_529
timestamp 1636968456
transform 1 0 50692 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_541
timestamp 1636968456
transform 1 0 51796 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_553
timestamp 1
transform 1 0 52900 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_559
timestamp 1
transform 1 0 53452 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_561
timestamp 1636968456
transform 1 0 53636 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_573
timestamp 1636968456
transform 1 0 54740 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_585
timestamp 1636968456
transform 1 0 55844 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_597
timestamp 1636968456
transform 1 0 56948 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_609
timestamp 1
transform 1 0 58052 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_615
timestamp 1
transform 1 0 58604 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_617
timestamp 1636968456
transform 1 0 58788 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_629
timestamp 1636968456
transform 1 0 59892 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_641
timestamp 1636968456
transform 1 0 60996 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_653
timestamp 1636968456
transform 1 0 62100 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_665
timestamp 1
transform 1 0 63204 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_671
timestamp 1
transform 1 0 63756 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_673
timestamp 1636968456
transform 1 0 63940 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_685
timestamp 1636968456
transform 1 0 65044 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_697
timestamp 1636968456
transform 1 0 66148 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_709
timestamp 1636968456
transform 1 0 67252 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_721
timestamp 1
transform 1 0 68356 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_727
timestamp 1
transform 1 0 68908 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_729
timestamp 1636968456
transform 1 0 69092 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_741
timestamp 1636968456
transform 1 0 70196 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_753
timestamp 1636968456
transform 1 0 71300 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_765
timestamp 1636968456
transform 1 0 72404 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_777
timestamp 1
transform 1 0 73508 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_783
timestamp 1
transform 1 0 74060 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_785
timestamp 1636968456
transform 1 0 74244 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_797
timestamp 1636968456
transform 1 0 75348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_809
timestamp 1636968456
transform 1 0 76452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_821
timestamp 1
transform 1 0 77556 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1636968456
transform 1 0 2300 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636968456
transform 1 0 3404 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1
transform 1 0 4508 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1636968456
transform 1 0 4692 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1636968456
transform 1 0 5796 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1636968456
transform 1 0 6900 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_65
timestamp 1636968456
transform 1 0 8004 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1
transform 1 0 9108 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1
transform 1 0 9660 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_85
timestamp 1636968456
transform 1 0 9844 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_97
timestamp 1636968456
transform 1 0 10948 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_109
timestamp 1636968456
transform 1 0 12052 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_121
timestamp 1636968456
transform 1 0 13156 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_133
timestamp 1
transform 1 0 14260 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1
transform 1 0 14812 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_141
timestamp 1636968456
transform 1 0 14996 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_153
timestamp 1636968456
transform 1 0 16100 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_165
timestamp 1636968456
transform 1 0 17204 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_177
timestamp 1636968456
transform 1 0 18308 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_189
timestamp 1
transform 1 0 19412 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_195
timestamp 1
transform 1 0 19964 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_197
timestamp 1636968456
transform 1 0 20148 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_209
timestamp 1636968456
transform 1 0 21252 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_221
timestamp 1636968456
transform 1 0 22356 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_233
timestamp 1636968456
transform 1 0 23460 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_245
timestamp 1
transform 1 0 24564 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_251
timestamp 1
transform 1 0 25116 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_253
timestamp 1636968456
transform 1 0 25300 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_265
timestamp 1636968456
transform 1 0 26404 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_277
timestamp 1636968456
transform 1 0 27508 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_289
timestamp 1636968456
transform 1 0 28612 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_301
timestamp 1
transform 1 0 29716 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_307
timestamp 1
transform 1 0 30268 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_309
timestamp 1636968456
transform 1 0 30452 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_321
timestamp 1636968456
transform 1 0 31556 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_333
timestamp 1636968456
transform 1 0 32660 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_345
timestamp 1636968456
transform 1 0 33764 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_357
timestamp 1
transform 1 0 34868 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_363
timestamp 1
transform 1 0 35420 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_365
timestamp 1636968456
transform 1 0 35604 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_377
timestamp 1636968456
transform 1 0 36708 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_389
timestamp 1636968456
transform 1 0 37812 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_401
timestamp 1636968456
transform 1 0 38916 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_413
timestamp 1
transform 1 0 40020 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_419
timestamp 1
transform 1 0 40572 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_421
timestamp 1636968456
transform 1 0 40756 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_433
timestamp 1636968456
transform 1 0 41860 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_445
timestamp 1636968456
transform 1 0 42964 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_457
timestamp 1636968456
transform 1 0 44068 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_469
timestamp 1
transform 1 0 45172 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_475
timestamp 1
transform 1 0 45724 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_477
timestamp 1636968456
transform 1 0 45908 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_489
timestamp 1636968456
transform 1 0 47012 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_501
timestamp 1636968456
transform 1 0 48116 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_513
timestamp 1636968456
transform 1 0 49220 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_525
timestamp 1
transform 1 0 50324 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1
transform 1 0 50876 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_533
timestamp 1636968456
transform 1 0 51060 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_545
timestamp 1636968456
transform 1 0 52164 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_557
timestamp 1636968456
transform 1 0 53268 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_569
timestamp 1636968456
transform 1 0 54372 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_581
timestamp 1
transform 1 0 55476 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_587
timestamp 1
transform 1 0 56028 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_589
timestamp 1636968456
transform 1 0 56212 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_601
timestamp 1636968456
transform 1 0 57316 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_613
timestamp 1636968456
transform 1 0 58420 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_625
timestamp 1636968456
transform 1 0 59524 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_637
timestamp 1
transform 1 0 60628 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_643
timestamp 1
transform 1 0 61180 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_645
timestamp 1636968456
transform 1 0 61364 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_657
timestamp 1636968456
transform 1 0 62468 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_669
timestamp 1636968456
transform 1 0 63572 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_681
timestamp 1636968456
transform 1 0 64676 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_693
timestamp 1
transform 1 0 65780 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_699
timestamp 1
transform 1 0 66332 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_701
timestamp 1636968456
transform 1 0 66516 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_713
timestamp 1636968456
transform 1 0 67620 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_725
timestamp 1636968456
transform 1 0 68724 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_737
timestamp 1636968456
transform 1 0 69828 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_749
timestamp 1
transform 1 0 70932 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_755
timestamp 1
transform 1 0 71484 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_757
timestamp 1636968456
transform 1 0 71668 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_769
timestamp 1636968456
transform 1 0 72772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_781
timestamp 1636968456
transform 1 0 73876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_793
timestamp 1636968456
transform 1 0 74980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_805
timestamp 1
transform 1 0 76084 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_811
timestamp 1
transform 1 0 76636 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_813
timestamp 1
transform 1 0 76820 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_821
timestamp 1
transform 1 0 77556 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1636968456
transform 1 0 2300 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1636968456
transform 1 0 3404 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_27
timestamp 1636968456
transform 1 0 4508 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_39
timestamp 1636968456
transform 1 0 5612 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_51
timestamp 1
transform 1 0 6716 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1
transform 1 0 7084 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1636968456
transform 1 0 7268 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_69
timestamp 1636968456
transform 1 0 8372 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_81
timestamp 1636968456
transform 1 0 9476 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_93
timestamp 1636968456
transform 1 0 10580 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_105
timestamp 1
transform 1 0 11684 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_111
timestamp 1
transform 1 0 12236 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_113
timestamp 1636968456
transform 1 0 12420 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_125
timestamp 1636968456
transform 1 0 13524 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_137
timestamp 1636968456
transform 1 0 14628 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_149
timestamp 1636968456
transform 1 0 15732 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_161
timestamp 1
transform 1 0 16836 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_167
timestamp 1
transform 1 0 17388 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_169
timestamp 1636968456
transform 1 0 17572 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_181
timestamp 1636968456
transform 1 0 18676 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_193
timestamp 1636968456
transform 1 0 19780 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_205
timestamp 1636968456
transform 1 0 20884 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_217
timestamp 1
transform 1 0 21988 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_223
timestamp 1
transform 1 0 22540 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_225
timestamp 1636968456
transform 1 0 22724 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_237
timestamp 1636968456
transform 1 0 23828 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_249
timestamp 1636968456
transform 1 0 24932 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_261
timestamp 1636968456
transform 1 0 26036 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_273
timestamp 1
transform 1 0 27140 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_279
timestamp 1
transform 1 0 27692 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_281
timestamp 1636968456
transform 1 0 27876 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_293
timestamp 1636968456
transform 1 0 28980 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_305
timestamp 1636968456
transform 1 0 30084 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_317
timestamp 1636968456
transform 1 0 31188 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_329
timestamp 1
transform 1 0 32292 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_335
timestamp 1
transform 1 0 32844 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_337
timestamp 1636968456
transform 1 0 33028 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_349
timestamp 1636968456
transform 1 0 34132 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_361
timestamp 1636968456
transform 1 0 35236 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_373
timestamp 1636968456
transform 1 0 36340 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_385
timestamp 1
transform 1 0 37444 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_391
timestamp 1
transform 1 0 37996 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_393
timestamp 1636968456
transform 1 0 38180 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_405
timestamp 1636968456
transform 1 0 39284 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_417
timestamp 1636968456
transform 1 0 40388 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_429
timestamp 1636968456
transform 1 0 41492 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_441
timestamp 1
transform 1 0 42596 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_447
timestamp 1
transform 1 0 43148 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_449
timestamp 1636968456
transform 1 0 43332 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_461
timestamp 1636968456
transform 1 0 44436 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_473
timestamp 1636968456
transform 1 0 45540 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_485
timestamp 1636968456
transform 1 0 46644 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_497
timestamp 1
transform 1 0 47748 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_503
timestamp 1
transform 1 0 48300 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_505
timestamp 1636968456
transform 1 0 48484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_517
timestamp 1636968456
transform 1 0 49588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_529
timestamp 1636968456
transform 1 0 50692 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_541
timestamp 1636968456
transform 1 0 51796 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_553
timestamp 1
transform 1 0 52900 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_559
timestamp 1
transform 1 0 53452 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_561
timestamp 1636968456
transform 1 0 53636 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_573
timestamp 1636968456
transform 1 0 54740 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_585
timestamp 1636968456
transform 1 0 55844 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_597
timestamp 1636968456
transform 1 0 56948 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_609
timestamp 1
transform 1 0 58052 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_615
timestamp 1
transform 1 0 58604 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_617
timestamp 1636968456
transform 1 0 58788 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_629
timestamp 1636968456
transform 1 0 59892 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_641
timestamp 1636968456
transform 1 0 60996 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_653
timestamp 1636968456
transform 1 0 62100 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_665
timestamp 1
transform 1 0 63204 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_671
timestamp 1
transform 1 0 63756 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_673
timestamp 1636968456
transform 1 0 63940 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_685
timestamp 1636968456
transform 1 0 65044 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_697
timestamp 1636968456
transform 1 0 66148 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_709
timestamp 1636968456
transform 1 0 67252 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_721
timestamp 1
transform 1 0 68356 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_727
timestamp 1
transform 1 0 68908 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_729
timestamp 1636968456
transform 1 0 69092 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_741
timestamp 1636968456
transform 1 0 70196 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_753
timestamp 1636968456
transform 1 0 71300 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_765
timestamp 1636968456
transform 1 0 72404 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_777
timestamp 1
transform 1 0 73508 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_783
timestamp 1
transform 1 0 74060 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_785
timestamp 1636968456
transform 1 0 74244 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_797
timestamp 1636968456
transform 1 0 75348 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_809
timestamp 1636968456
transform 1 0 76452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_821
timestamp 1
transform 1 0 77556 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1636968456
transform 1 0 2300 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1636968456
transform 1 0 3404 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1
transform 1 0 4508 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1636968456
transform 1 0 4692 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_41
timestamp 1636968456
transform 1 0 5796 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_53
timestamp 1636968456
transform 1 0 6900 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_65
timestamp 1636968456
transform 1 0 8004 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1
transform 1 0 9108 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1
transform 1 0 9660 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_85
timestamp 1636968456
transform 1 0 9844 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_97
timestamp 1636968456
transform 1 0 10948 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_109
timestamp 1636968456
transform 1 0 12052 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_121
timestamp 1636968456
transform 1 0 13156 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_133
timestamp 1
transform 1 0 14260 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_139
timestamp 1
transform 1 0 14812 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_141
timestamp 1636968456
transform 1 0 14996 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_153
timestamp 1636968456
transform 1 0 16100 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_165
timestamp 1636968456
transform 1 0 17204 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_177
timestamp 1636968456
transform 1 0 18308 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_189
timestamp 1
transform 1 0 19412 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_195
timestamp 1
transform 1 0 19964 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_197
timestamp 1636968456
transform 1 0 20148 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_209
timestamp 1636968456
transform 1 0 21252 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_221
timestamp 1636968456
transform 1 0 22356 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_233
timestamp 1636968456
transform 1 0 23460 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_245
timestamp 1
transform 1 0 24564 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_251
timestamp 1
transform 1 0 25116 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_253
timestamp 1636968456
transform 1 0 25300 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_265
timestamp 1636968456
transform 1 0 26404 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_277
timestamp 1636968456
transform 1 0 27508 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_289
timestamp 1636968456
transform 1 0 28612 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_301
timestamp 1
transform 1 0 29716 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_307
timestamp 1
transform 1 0 30268 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_309
timestamp 1636968456
transform 1 0 30452 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_321
timestamp 1636968456
transform 1 0 31556 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_333
timestamp 1636968456
transform 1 0 32660 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_345
timestamp 1636968456
transform 1 0 33764 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_357
timestamp 1
transform 1 0 34868 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_363
timestamp 1
transform 1 0 35420 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_365
timestamp 1636968456
transform 1 0 35604 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_377
timestamp 1636968456
transform 1 0 36708 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_389
timestamp 1636968456
transform 1 0 37812 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_401
timestamp 1636968456
transform 1 0 38916 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_413
timestamp 1
transform 1 0 40020 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_419
timestamp 1
transform 1 0 40572 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_421
timestamp 1636968456
transform 1 0 40756 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_433
timestamp 1636968456
transform 1 0 41860 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_445
timestamp 1636968456
transform 1 0 42964 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_457
timestamp 1636968456
transform 1 0 44068 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_469
timestamp 1
transform 1 0 45172 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_475
timestamp 1
transform 1 0 45724 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_477
timestamp 1636968456
transform 1 0 45908 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_489
timestamp 1636968456
transform 1 0 47012 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_501
timestamp 1636968456
transform 1 0 48116 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_513
timestamp 1636968456
transform 1 0 49220 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_525
timestamp 1
transform 1 0 50324 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1
transform 1 0 50876 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_533
timestamp 1636968456
transform 1 0 51060 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_545
timestamp 1636968456
transform 1 0 52164 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_557
timestamp 1636968456
transform 1 0 53268 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_569
timestamp 1636968456
transform 1 0 54372 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_581
timestamp 1
transform 1 0 55476 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_587
timestamp 1
transform 1 0 56028 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_589
timestamp 1636968456
transform 1 0 56212 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_601
timestamp 1636968456
transform 1 0 57316 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_613
timestamp 1636968456
transform 1 0 58420 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_625
timestamp 1636968456
transform 1 0 59524 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_637
timestamp 1
transform 1 0 60628 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_643
timestamp 1
transform 1 0 61180 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_645
timestamp 1636968456
transform 1 0 61364 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_657
timestamp 1636968456
transform 1 0 62468 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_669
timestamp 1636968456
transform 1 0 63572 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_681
timestamp 1636968456
transform 1 0 64676 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_693
timestamp 1
transform 1 0 65780 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_699
timestamp 1
transform 1 0 66332 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_701
timestamp 1636968456
transform 1 0 66516 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_713
timestamp 1636968456
transform 1 0 67620 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_725
timestamp 1636968456
transform 1 0 68724 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_737
timestamp 1636968456
transform 1 0 69828 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_749
timestamp 1
transform 1 0 70932 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_755
timestamp 1
transform 1 0 71484 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_757
timestamp 1636968456
transform 1 0 71668 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_769
timestamp 1636968456
transform 1 0 72772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_781
timestamp 1636968456
transform 1 0 73876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_793
timestamp 1636968456
transform 1 0 74980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_805
timestamp 1
transform 1 0 76084 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_811
timestamp 1
transform 1 0 76636 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_813
timestamp 1
transform 1 0 76820 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_821
timestamp 1
transform 1 0 77556 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_3
timestamp 1636968456
transform 1 0 2300 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_15
timestamp 1636968456
transform 1 0 3404 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_27
timestamp 1636968456
transform 1 0 4508 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_39
timestamp 1636968456
transform 1 0 5612 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1
transform 1 0 6716 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1
transform 1 0 7084 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_57
timestamp 1636968456
transform 1 0 7268 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_69
timestamp 1636968456
transform 1 0 8372 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_81
timestamp 1636968456
transform 1 0 9476 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_93
timestamp 1636968456
transform 1 0 10580 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_105
timestamp 1
transform 1 0 11684 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_111
timestamp 1
transform 1 0 12236 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_113
timestamp 1636968456
transform 1 0 12420 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_125
timestamp 1636968456
transform 1 0 13524 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_137
timestamp 1636968456
transform 1 0 14628 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_149
timestamp 1636968456
transform 1 0 15732 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_161
timestamp 1
transform 1 0 16836 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_167
timestamp 1
transform 1 0 17388 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_169
timestamp 1636968456
transform 1 0 17572 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_181
timestamp 1636968456
transform 1 0 18676 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_193
timestamp 1636968456
transform 1 0 19780 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_205
timestamp 1636968456
transform 1 0 20884 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_217
timestamp 1
transform 1 0 21988 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_223
timestamp 1
transform 1 0 22540 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_225
timestamp 1636968456
transform 1 0 22724 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_237
timestamp 1636968456
transform 1 0 23828 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_249
timestamp 1636968456
transform 1 0 24932 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_261
timestamp 1636968456
transform 1 0 26036 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_273
timestamp 1
transform 1 0 27140 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_279
timestamp 1
transform 1 0 27692 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_281
timestamp 1636968456
transform 1 0 27876 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_293
timestamp 1636968456
transform 1 0 28980 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_305
timestamp 1636968456
transform 1 0 30084 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_317
timestamp 1636968456
transform 1 0 31188 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_329
timestamp 1
transform 1 0 32292 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_335
timestamp 1
transform 1 0 32844 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_337
timestamp 1636968456
transform 1 0 33028 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_349
timestamp 1636968456
transform 1 0 34132 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_361
timestamp 1636968456
transform 1 0 35236 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_373
timestamp 1636968456
transform 1 0 36340 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_385
timestamp 1
transform 1 0 37444 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_391
timestamp 1
transform 1 0 37996 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_393
timestamp 1636968456
transform 1 0 38180 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_405
timestamp 1636968456
transform 1 0 39284 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_417
timestamp 1636968456
transform 1 0 40388 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_429
timestamp 1636968456
transform 1 0 41492 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_441
timestamp 1
transform 1 0 42596 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_447
timestamp 1
transform 1 0 43148 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_449
timestamp 1636968456
transform 1 0 43332 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_461
timestamp 1636968456
transform 1 0 44436 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_473
timestamp 1636968456
transform 1 0 45540 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_485
timestamp 1636968456
transform 1 0 46644 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_497
timestamp 1
transform 1 0 47748 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_503
timestamp 1
transform 1 0 48300 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_505
timestamp 1636968456
transform 1 0 48484 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_517
timestamp 1636968456
transform 1 0 49588 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_529
timestamp 1636968456
transform 1 0 50692 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_541
timestamp 1636968456
transform 1 0 51796 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_553
timestamp 1
transform 1 0 52900 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_559
timestamp 1
transform 1 0 53452 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_561
timestamp 1636968456
transform 1 0 53636 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_573
timestamp 1636968456
transform 1 0 54740 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_585
timestamp 1636968456
transform 1 0 55844 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_597
timestamp 1636968456
transform 1 0 56948 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_609
timestamp 1
transform 1 0 58052 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_615
timestamp 1
transform 1 0 58604 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_617
timestamp 1636968456
transform 1 0 58788 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_629
timestamp 1636968456
transform 1 0 59892 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_641
timestamp 1636968456
transform 1 0 60996 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_653
timestamp 1636968456
transform 1 0 62100 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_665
timestamp 1
transform 1 0 63204 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_671
timestamp 1
transform 1 0 63756 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_673
timestamp 1636968456
transform 1 0 63940 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_685
timestamp 1636968456
transform 1 0 65044 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_697
timestamp 1636968456
transform 1 0 66148 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_709
timestamp 1636968456
transform 1 0 67252 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_721
timestamp 1
transform 1 0 68356 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_727
timestamp 1
transform 1 0 68908 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_729
timestamp 1636968456
transform 1 0 69092 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_741
timestamp 1636968456
transform 1 0 70196 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_753
timestamp 1636968456
transform 1 0 71300 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_765
timestamp 1636968456
transform 1 0 72404 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_777
timestamp 1
transform 1 0 73508 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_783
timestamp 1
transform 1 0 74060 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_785
timestamp 1636968456
transform 1 0 74244 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_797
timestamp 1636968456
transform 1 0 75348 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_809
timestamp 1636968456
transform 1 0 76452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_109_821
timestamp 1
transform 1 0 77556 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_3
timestamp 1636968456
transform 1 0 2300 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_15
timestamp 1636968456
transform 1 0 3404 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1
transform 1 0 4508 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1636968456
transform 1 0 4692 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_41
timestamp 1636968456
transform 1 0 5796 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_53
timestamp 1636968456
transform 1 0 6900 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_65
timestamp 1636968456
transform 1 0 8004 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1
transform 1 0 9108 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1
transform 1 0 9660 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_85
timestamp 1636968456
transform 1 0 9844 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_97
timestamp 1636968456
transform 1 0 10948 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_109
timestamp 1636968456
transform 1 0 12052 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_121
timestamp 1636968456
transform 1 0 13156 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_133
timestamp 1
transform 1 0 14260 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_139
timestamp 1
transform 1 0 14812 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_141
timestamp 1636968456
transform 1 0 14996 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_153
timestamp 1636968456
transform 1 0 16100 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_165
timestamp 1636968456
transform 1 0 17204 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_177
timestamp 1636968456
transform 1 0 18308 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_189
timestamp 1
transform 1 0 19412 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_195
timestamp 1
transform 1 0 19964 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_197
timestamp 1636968456
transform 1 0 20148 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_209
timestamp 1636968456
transform 1 0 21252 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_221
timestamp 1636968456
transform 1 0 22356 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_233
timestamp 1636968456
transform 1 0 23460 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_245
timestamp 1
transform 1 0 24564 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_251
timestamp 1
transform 1 0 25116 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_253
timestamp 1636968456
transform 1 0 25300 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_265
timestamp 1636968456
transform 1 0 26404 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_277
timestamp 1636968456
transform 1 0 27508 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_289
timestamp 1636968456
transform 1 0 28612 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_301
timestamp 1
transform 1 0 29716 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_307
timestamp 1
transform 1 0 30268 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_309
timestamp 1636968456
transform 1 0 30452 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_321
timestamp 1636968456
transform 1 0 31556 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_333
timestamp 1636968456
transform 1 0 32660 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_345
timestamp 1636968456
transform 1 0 33764 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_357
timestamp 1
transform 1 0 34868 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_363
timestamp 1
transform 1 0 35420 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_365
timestamp 1636968456
transform 1 0 35604 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_377
timestamp 1636968456
transform 1 0 36708 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_389
timestamp 1636968456
transform 1 0 37812 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_401
timestamp 1636968456
transform 1 0 38916 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_413
timestamp 1
transform 1 0 40020 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_419
timestamp 1
transform 1 0 40572 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_421
timestamp 1636968456
transform 1 0 40756 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_433
timestamp 1636968456
transform 1 0 41860 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_445
timestamp 1636968456
transform 1 0 42964 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_457
timestamp 1636968456
transform 1 0 44068 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_469
timestamp 1
transform 1 0 45172 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_475
timestamp 1
transform 1 0 45724 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_477
timestamp 1636968456
transform 1 0 45908 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_489
timestamp 1636968456
transform 1 0 47012 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_501
timestamp 1636968456
transform 1 0 48116 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_513
timestamp 1636968456
transform 1 0 49220 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_525
timestamp 1
transform 1 0 50324 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_531
timestamp 1
transform 1 0 50876 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_533
timestamp 1636968456
transform 1 0 51060 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_545
timestamp 1636968456
transform 1 0 52164 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_557
timestamp 1636968456
transform 1 0 53268 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_569
timestamp 1636968456
transform 1 0 54372 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_581
timestamp 1
transform 1 0 55476 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_587
timestamp 1
transform 1 0 56028 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_589
timestamp 1636968456
transform 1 0 56212 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_601
timestamp 1636968456
transform 1 0 57316 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_613
timestamp 1636968456
transform 1 0 58420 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_625
timestamp 1636968456
transform 1 0 59524 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_637
timestamp 1
transform 1 0 60628 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_643
timestamp 1
transform 1 0 61180 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_645
timestamp 1636968456
transform 1 0 61364 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_657
timestamp 1636968456
transform 1 0 62468 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_669
timestamp 1636968456
transform 1 0 63572 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_681
timestamp 1636968456
transform 1 0 64676 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_693
timestamp 1
transform 1 0 65780 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_699
timestamp 1
transform 1 0 66332 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_701
timestamp 1636968456
transform 1 0 66516 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_713
timestamp 1636968456
transform 1 0 67620 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_725
timestamp 1636968456
transform 1 0 68724 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_737
timestamp 1636968456
transform 1 0 69828 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_749
timestamp 1
transform 1 0 70932 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_755
timestamp 1
transform 1 0 71484 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_757
timestamp 1636968456
transform 1 0 71668 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_769
timestamp 1636968456
transform 1 0 72772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_781
timestamp 1636968456
transform 1 0 73876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_793
timestamp 1636968456
transform 1 0 74980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_805
timestamp 1
transform 1 0 76084 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_811
timestamp 1
transform 1 0 76636 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_813
timestamp 1
transform 1 0 76820 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_110_821
timestamp 1
transform 1 0 77556 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1636968456
transform 1 0 2300 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1636968456
transform 1 0 3404 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_27
timestamp 1636968456
transform 1 0 4508 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_39
timestamp 1636968456
transform 1 0 5612 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1
transform 1 0 6716 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1
transform 1 0 7084 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_57
timestamp 1636968456
transform 1 0 7268 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_69
timestamp 1636968456
transform 1 0 8372 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_81
timestamp 1636968456
transform 1 0 9476 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_93
timestamp 1636968456
transform 1 0 10580 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_105
timestamp 1
transform 1 0 11684 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_111
timestamp 1
transform 1 0 12236 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_113
timestamp 1636968456
transform 1 0 12420 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_125
timestamp 1636968456
transform 1 0 13524 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_137
timestamp 1636968456
transform 1 0 14628 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_149
timestamp 1636968456
transform 1 0 15732 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_161
timestamp 1
transform 1 0 16836 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_167
timestamp 1
transform 1 0 17388 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_169
timestamp 1636968456
transform 1 0 17572 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_181
timestamp 1636968456
transform 1 0 18676 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_193
timestamp 1636968456
transform 1 0 19780 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_205
timestamp 1636968456
transform 1 0 20884 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_217
timestamp 1
transform 1 0 21988 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_223
timestamp 1
transform 1 0 22540 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_225
timestamp 1636968456
transform 1 0 22724 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_237
timestamp 1636968456
transform 1 0 23828 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_249
timestamp 1636968456
transform 1 0 24932 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_261
timestamp 1636968456
transform 1 0 26036 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_273
timestamp 1
transform 1 0 27140 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_279
timestamp 1
transform 1 0 27692 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_281
timestamp 1636968456
transform 1 0 27876 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_293
timestamp 1636968456
transform 1 0 28980 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_305
timestamp 1636968456
transform 1 0 30084 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_317
timestamp 1636968456
transform 1 0 31188 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_329
timestamp 1
transform 1 0 32292 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_335
timestamp 1
transform 1 0 32844 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_337
timestamp 1636968456
transform 1 0 33028 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_349
timestamp 1636968456
transform 1 0 34132 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_361
timestamp 1636968456
transform 1 0 35236 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_373
timestamp 1636968456
transform 1 0 36340 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_385
timestamp 1
transform 1 0 37444 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_391
timestamp 1
transform 1 0 37996 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_393
timestamp 1636968456
transform 1 0 38180 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_405
timestamp 1636968456
transform 1 0 39284 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_417
timestamp 1636968456
transform 1 0 40388 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_429
timestamp 1636968456
transform 1 0 41492 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_441
timestamp 1
transform 1 0 42596 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_447
timestamp 1
transform 1 0 43148 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_449
timestamp 1636968456
transform 1 0 43332 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_461
timestamp 1636968456
transform 1 0 44436 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_473
timestamp 1636968456
transform 1 0 45540 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_485
timestamp 1636968456
transform 1 0 46644 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_497
timestamp 1
transform 1 0 47748 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_503
timestamp 1
transform 1 0 48300 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_505
timestamp 1636968456
transform 1 0 48484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_517
timestamp 1636968456
transform 1 0 49588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_529
timestamp 1636968456
transform 1 0 50692 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_541
timestamp 1636968456
transform 1 0 51796 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_553
timestamp 1
transform 1 0 52900 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_559
timestamp 1
transform 1 0 53452 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_561
timestamp 1636968456
transform 1 0 53636 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_573
timestamp 1636968456
transform 1 0 54740 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_585
timestamp 1636968456
transform 1 0 55844 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_597
timestamp 1636968456
transform 1 0 56948 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_609
timestamp 1
transform 1 0 58052 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_615
timestamp 1
transform 1 0 58604 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_617
timestamp 1636968456
transform 1 0 58788 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_629
timestamp 1636968456
transform 1 0 59892 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_641
timestamp 1636968456
transform 1 0 60996 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_653
timestamp 1636968456
transform 1 0 62100 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_665
timestamp 1
transform 1 0 63204 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_671
timestamp 1
transform 1 0 63756 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_673
timestamp 1636968456
transform 1 0 63940 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_685
timestamp 1636968456
transform 1 0 65044 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_697
timestamp 1636968456
transform 1 0 66148 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_709
timestamp 1636968456
transform 1 0 67252 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_721
timestamp 1
transform 1 0 68356 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_727
timestamp 1
transform 1 0 68908 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_729
timestamp 1636968456
transform 1 0 69092 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_741
timestamp 1636968456
transform 1 0 70196 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_753
timestamp 1636968456
transform 1 0 71300 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_765
timestamp 1636968456
transform 1 0 72404 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_777
timestamp 1
transform 1 0 73508 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_783
timestamp 1
transform 1 0 74060 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_785
timestamp 1636968456
transform 1 0 74244 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_797
timestamp 1636968456
transform 1 0 75348 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_809
timestamp 1636968456
transform 1 0 76452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_111_821
timestamp 1
transform 1 0 77556 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_3
timestamp 1636968456
transform 1 0 2300 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_15
timestamp 1636968456
transform 1 0 3404 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1
transform 1 0 4508 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1636968456
transform 1 0 4692 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_41
timestamp 1636968456
transform 1 0 5796 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_53
timestamp 1636968456
transform 1 0 6900 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_65
timestamp 1636968456
transform 1 0 8004 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1
transform 1 0 9108 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1
transform 1 0 9660 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_85
timestamp 1636968456
transform 1 0 9844 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_97
timestamp 1636968456
transform 1 0 10948 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_109
timestamp 1636968456
transform 1 0 12052 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_121
timestamp 1636968456
transform 1 0 13156 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_133
timestamp 1
transform 1 0 14260 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_139
timestamp 1
transform 1 0 14812 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_141
timestamp 1636968456
transform 1 0 14996 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_153
timestamp 1636968456
transform 1 0 16100 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_165
timestamp 1636968456
transform 1 0 17204 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_177
timestamp 1636968456
transform 1 0 18308 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_189
timestamp 1
transform 1 0 19412 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_195
timestamp 1
transform 1 0 19964 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_197
timestamp 1636968456
transform 1 0 20148 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_209
timestamp 1636968456
transform 1 0 21252 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_221
timestamp 1636968456
transform 1 0 22356 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_233
timestamp 1636968456
transform 1 0 23460 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_245
timestamp 1
transform 1 0 24564 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_251
timestamp 1
transform 1 0 25116 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_253
timestamp 1636968456
transform 1 0 25300 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_265
timestamp 1636968456
transform 1 0 26404 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_277
timestamp 1636968456
transform 1 0 27508 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_289
timestamp 1636968456
transform 1 0 28612 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_301
timestamp 1
transform 1 0 29716 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_307
timestamp 1
transform 1 0 30268 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_309
timestamp 1636968456
transform 1 0 30452 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_321
timestamp 1636968456
transform 1 0 31556 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_333
timestamp 1636968456
transform 1 0 32660 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_345
timestamp 1636968456
transform 1 0 33764 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_357
timestamp 1
transform 1 0 34868 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_363
timestamp 1
transform 1 0 35420 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_365
timestamp 1636968456
transform 1 0 35604 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_377
timestamp 1636968456
transform 1 0 36708 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_389
timestamp 1636968456
transform 1 0 37812 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_401
timestamp 1636968456
transform 1 0 38916 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_413
timestamp 1
transform 1 0 40020 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_419
timestamp 1
transform 1 0 40572 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_421
timestamp 1636968456
transform 1 0 40756 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_433
timestamp 1636968456
transform 1 0 41860 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_445
timestamp 1636968456
transform 1 0 42964 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_457
timestamp 1636968456
transform 1 0 44068 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_469
timestamp 1
transform 1 0 45172 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_475
timestamp 1
transform 1 0 45724 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_477
timestamp 1636968456
transform 1 0 45908 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_489
timestamp 1636968456
transform 1 0 47012 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_501
timestamp 1636968456
transform 1 0 48116 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_513
timestamp 1636968456
transform 1 0 49220 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_525
timestamp 1
transform 1 0 50324 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_531
timestamp 1
transform 1 0 50876 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_533
timestamp 1636968456
transform 1 0 51060 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_545
timestamp 1636968456
transform 1 0 52164 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_557
timestamp 1636968456
transform 1 0 53268 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_569
timestamp 1636968456
transform 1 0 54372 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_581
timestamp 1
transform 1 0 55476 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_587
timestamp 1
transform 1 0 56028 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_589
timestamp 1636968456
transform 1 0 56212 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_601
timestamp 1636968456
transform 1 0 57316 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_613
timestamp 1636968456
transform 1 0 58420 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_625
timestamp 1636968456
transform 1 0 59524 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_637
timestamp 1
transform 1 0 60628 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_643
timestamp 1
transform 1 0 61180 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_645
timestamp 1636968456
transform 1 0 61364 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_657
timestamp 1636968456
transform 1 0 62468 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_669
timestamp 1636968456
transform 1 0 63572 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_681
timestamp 1636968456
transform 1 0 64676 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_693
timestamp 1
transform 1 0 65780 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_699
timestamp 1
transform 1 0 66332 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_701
timestamp 1636968456
transform 1 0 66516 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_713
timestamp 1636968456
transform 1 0 67620 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_725
timestamp 1636968456
transform 1 0 68724 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_737
timestamp 1636968456
transform 1 0 69828 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_749
timestamp 1
transform 1 0 70932 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_755
timestamp 1
transform 1 0 71484 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_757
timestamp 1636968456
transform 1 0 71668 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_769
timestamp 1636968456
transform 1 0 72772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_781
timestamp 1636968456
transform 1 0 73876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_793
timestamp 1636968456
transform 1 0 74980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_805
timestamp 1
transform 1 0 76084 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_811
timestamp 1
transform 1 0 76636 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_813
timestamp 1
transform 1 0 76820 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_112_821
timestamp 1
transform 1 0 77556 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636968456
transform 1 0 2300 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636968456
transform 1 0 3404 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1636968456
transform 1 0 4508 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_39
timestamp 1636968456
transform 1 0 5612 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1
transform 1 0 6716 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1
transform 1 0 7084 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_57
timestamp 1636968456
transform 1 0 7268 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_69
timestamp 1636968456
transform 1 0 8372 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_81
timestamp 1636968456
transform 1 0 9476 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_93
timestamp 1636968456
transform 1 0 10580 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_105
timestamp 1
transform 1 0 11684 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_111
timestamp 1
transform 1 0 12236 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_113
timestamp 1636968456
transform 1 0 12420 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_125
timestamp 1636968456
transform 1 0 13524 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_137
timestamp 1636968456
transform 1 0 14628 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_149
timestamp 1636968456
transform 1 0 15732 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_161
timestamp 1
transform 1 0 16836 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_167
timestamp 1
transform 1 0 17388 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_169
timestamp 1636968456
transform 1 0 17572 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_181
timestamp 1636968456
transform 1 0 18676 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_193
timestamp 1636968456
transform 1 0 19780 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_205
timestamp 1636968456
transform 1 0 20884 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_217
timestamp 1
transform 1 0 21988 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_223
timestamp 1
transform 1 0 22540 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_225
timestamp 1636968456
transform 1 0 22724 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_237
timestamp 1636968456
transform 1 0 23828 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_249
timestamp 1636968456
transform 1 0 24932 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_261
timestamp 1636968456
transform 1 0 26036 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_273
timestamp 1
transform 1 0 27140 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_279
timestamp 1
transform 1 0 27692 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_281
timestamp 1636968456
transform 1 0 27876 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_293
timestamp 1636968456
transform 1 0 28980 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_305
timestamp 1636968456
transform 1 0 30084 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_317
timestamp 1636968456
transform 1 0 31188 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_329
timestamp 1
transform 1 0 32292 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_335
timestamp 1
transform 1 0 32844 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_337
timestamp 1636968456
transform 1 0 33028 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_349
timestamp 1636968456
transform 1 0 34132 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_361
timestamp 1636968456
transform 1 0 35236 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_373
timestamp 1636968456
transform 1 0 36340 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_385
timestamp 1
transform 1 0 37444 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_391
timestamp 1
transform 1 0 37996 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_393
timestamp 1636968456
transform 1 0 38180 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_405
timestamp 1636968456
transform 1 0 39284 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_417
timestamp 1636968456
transform 1 0 40388 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_429
timestamp 1636968456
transform 1 0 41492 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_441
timestamp 1
transform 1 0 42596 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_447
timestamp 1
transform 1 0 43148 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_449
timestamp 1636968456
transform 1 0 43332 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_461
timestamp 1636968456
transform 1 0 44436 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_473
timestamp 1636968456
transform 1 0 45540 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_485
timestamp 1636968456
transform 1 0 46644 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_497
timestamp 1
transform 1 0 47748 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_503
timestamp 1
transform 1 0 48300 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_505
timestamp 1636968456
transform 1 0 48484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_517
timestamp 1636968456
transform 1 0 49588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_529
timestamp 1636968456
transform 1 0 50692 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_541
timestamp 1636968456
transform 1 0 51796 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_553
timestamp 1
transform 1 0 52900 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_559
timestamp 1
transform 1 0 53452 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_561
timestamp 1636968456
transform 1 0 53636 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_573
timestamp 1636968456
transform 1 0 54740 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_585
timestamp 1636968456
transform 1 0 55844 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_597
timestamp 1636968456
transform 1 0 56948 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_609
timestamp 1
transform 1 0 58052 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_615
timestamp 1
transform 1 0 58604 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_617
timestamp 1636968456
transform 1 0 58788 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_629
timestamp 1636968456
transform 1 0 59892 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_641
timestamp 1636968456
transform 1 0 60996 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_653
timestamp 1636968456
transform 1 0 62100 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_665
timestamp 1
transform 1 0 63204 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_671
timestamp 1
transform 1 0 63756 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_673
timestamp 1636968456
transform 1 0 63940 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_685
timestamp 1636968456
transform 1 0 65044 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_697
timestamp 1636968456
transform 1 0 66148 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_709
timestamp 1636968456
transform 1 0 67252 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_721
timestamp 1
transform 1 0 68356 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_727
timestamp 1
transform 1 0 68908 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_729
timestamp 1636968456
transform 1 0 69092 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_741
timestamp 1636968456
transform 1 0 70196 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_753
timestamp 1636968456
transform 1 0 71300 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_765
timestamp 1636968456
transform 1 0 72404 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_777
timestamp 1
transform 1 0 73508 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_783
timestamp 1
transform 1 0 74060 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_785
timestamp 1636968456
transform 1 0 74244 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_797
timestamp 1636968456
transform 1 0 75348 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_809
timestamp 1636968456
transform 1 0 76452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_113_821
timestamp 1
transform 1 0 77556 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_3
timestamp 1636968456
transform 1 0 2300 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_15
timestamp 1636968456
transform 1 0 3404 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1
transform 1 0 4508 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1636968456
transform 1 0 4692 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_41
timestamp 1636968456
transform 1 0 5796 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_53
timestamp 1636968456
transform 1 0 6900 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_65
timestamp 1636968456
transform 1 0 8004 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1
transform 1 0 9108 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1
transform 1 0 9660 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_85
timestamp 1636968456
transform 1 0 9844 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_97
timestamp 1636968456
transform 1 0 10948 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_109
timestamp 1636968456
transform 1 0 12052 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_121
timestamp 1636968456
transform 1 0 13156 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_133
timestamp 1
transform 1 0 14260 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_139
timestamp 1
transform 1 0 14812 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_141
timestamp 1636968456
transform 1 0 14996 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_153
timestamp 1636968456
transform 1 0 16100 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_165
timestamp 1636968456
transform 1 0 17204 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_177
timestamp 1636968456
transform 1 0 18308 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_189
timestamp 1
transform 1 0 19412 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_195
timestamp 1
transform 1 0 19964 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_197
timestamp 1636968456
transform 1 0 20148 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_209
timestamp 1636968456
transform 1 0 21252 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_221
timestamp 1636968456
transform 1 0 22356 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_233
timestamp 1636968456
transform 1 0 23460 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_245
timestamp 1
transform 1 0 24564 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_251
timestamp 1
transform 1 0 25116 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_253
timestamp 1636968456
transform 1 0 25300 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_265
timestamp 1636968456
transform 1 0 26404 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_277
timestamp 1636968456
transform 1 0 27508 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_289
timestamp 1636968456
transform 1 0 28612 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_301
timestamp 1
transform 1 0 29716 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_307
timestamp 1
transform 1 0 30268 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_309
timestamp 1636968456
transform 1 0 30452 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_321
timestamp 1636968456
transform 1 0 31556 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_333
timestamp 1636968456
transform 1 0 32660 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_345
timestamp 1636968456
transform 1 0 33764 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_357
timestamp 1
transform 1 0 34868 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_363
timestamp 1
transform 1 0 35420 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_365
timestamp 1636968456
transform 1 0 35604 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_377
timestamp 1636968456
transform 1 0 36708 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_389
timestamp 1636968456
transform 1 0 37812 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_401
timestamp 1636968456
transform 1 0 38916 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_413
timestamp 1
transform 1 0 40020 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_419
timestamp 1
transform 1 0 40572 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_421
timestamp 1636968456
transform 1 0 40756 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_433
timestamp 1636968456
transform 1 0 41860 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_445
timestamp 1636968456
transform 1 0 42964 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_457
timestamp 1636968456
transform 1 0 44068 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_469
timestamp 1
transform 1 0 45172 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_475
timestamp 1
transform 1 0 45724 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_477
timestamp 1636968456
transform 1 0 45908 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_489
timestamp 1636968456
transform 1 0 47012 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_501
timestamp 1636968456
transform 1 0 48116 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_513
timestamp 1636968456
transform 1 0 49220 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_525
timestamp 1
transform 1 0 50324 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_531
timestamp 1
transform 1 0 50876 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_533
timestamp 1636968456
transform 1 0 51060 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_545
timestamp 1636968456
transform 1 0 52164 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_557
timestamp 1636968456
transform 1 0 53268 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_569
timestamp 1636968456
transform 1 0 54372 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_581
timestamp 1
transform 1 0 55476 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_587
timestamp 1
transform 1 0 56028 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_589
timestamp 1636968456
transform 1 0 56212 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_601
timestamp 1636968456
transform 1 0 57316 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_613
timestamp 1636968456
transform 1 0 58420 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_625
timestamp 1636968456
transform 1 0 59524 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_637
timestamp 1
transform 1 0 60628 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_643
timestamp 1
transform 1 0 61180 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_645
timestamp 1636968456
transform 1 0 61364 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_657
timestamp 1636968456
transform 1 0 62468 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_669
timestamp 1636968456
transform 1 0 63572 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_681
timestamp 1636968456
transform 1 0 64676 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_693
timestamp 1
transform 1 0 65780 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_699
timestamp 1
transform 1 0 66332 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_701
timestamp 1636968456
transform 1 0 66516 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_713
timestamp 1636968456
transform 1 0 67620 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_725
timestamp 1636968456
transform 1 0 68724 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_737
timestamp 1636968456
transform 1 0 69828 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_749
timestamp 1
transform 1 0 70932 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_755
timestamp 1
transform 1 0 71484 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_757
timestamp 1636968456
transform 1 0 71668 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_769
timestamp 1636968456
transform 1 0 72772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_781
timestamp 1636968456
transform 1 0 73876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_793
timestamp 1636968456
transform 1 0 74980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_805
timestamp 1
transform 1 0 76084 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_811
timestamp 1
transform 1 0 76636 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_813
timestamp 1
transform 1 0 76820 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_114_821
timestamp 1
transform 1 0 77556 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_3
timestamp 1636968456
transform 1 0 2300 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_15
timestamp 1636968456
transform 1 0 3404 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_27
timestamp 1636968456
transform 1 0 4508 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_39
timestamp 1636968456
transform 1 0 5612 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1
transform 1 0 6716 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1
transform 1 0 7084 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_57
timestamp 1636968456
transform 1 0 7268 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_69
timestamp 1636968456
transform 1 0 8372 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_81
timestamp 1636968456
transform 1 0 9476 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_93
timestamp 1636968456
transform 1 0 10580 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_105
timestamp 1
transform 1 0 11684 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_111
timestamp 1
transform 1 0 12236 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_113
timestamp 1636968456
transform 1 0 12420 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_125
timestamp 1636968456
transform 1 0 13524 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_137
timestamp 1636968456
transform 1 0 14628 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_149
timestamp 1636968456
transform 1 0 15732 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_161
timestamp 1
transform 1 0 16836 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_167
timestamp 1
transform 1 0 17388 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_169
timestamp 1636968456
transform 1 0 17572 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_181
timestamp 1636968456
transform 1 0 18676 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_193
timestamp 1636968456
transform 1 0 19780 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_205
timestamp 1636968456
transform 1 0 20884 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_217
timestamp 1
transform 1 0 21988 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_223
timestamp 1
transform 1 0 22540 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_225
timestamp 1636968456
transform 1 0 22724 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_237
timestamp 1636968456
transform 1 0 23828 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_249
timestamp 1636968456
transform 1 0 24932 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_261
timestamp 1636968456
transform 1 0 26036 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_273
timestamp 1
transform 1 0 27140 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_279
timestamp 1
transform 1 0 27692 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_281
timestamp 1636968456
transform 1 0 27876 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_293
timestamp 1636968456
transform 1 0 28980 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_305
timestamp 1636968456
transform 1 0 30084 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_317
timestamp 1636968456
transform 1 0 31188 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_329
timestamp 1
transform 1 0 32292 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_335
timestamp 1
transform 1 0 32844 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_337
timestamp 1636968456
transform 1 0 33028 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_349
timestamp 1636968456
transform 1 0 34132 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_361
timestamp 1636968456
transform 1 0 35236 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_373
timestamp 1636968456
transform 1 0 36340 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_385
timestamp 1
transform 1 0 37444 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_391
timestamp 1
transform 1 0 37996 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_393
timestamp 1636968456
transform 1 0 38180 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_405
timestamp 1636968456
transform 1 0 39284 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_417
timestamp 1636968456
transform 1 0 40388 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_429
timestamp 1636968456
transform 1 0 41492 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_441
timestamp 1
transform 1 0 42596 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_447
timestamp 1
transform 1 0 43148 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_449
timestamp 1636968456
transform 1 0 43332 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_461
timestamp 1636968456
transform 1 0 44436 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_473
timestamp 1636968456
transform 1 0 45540 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_485
timestamp 1636968456
transform 1 0 46644 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_497
timestamp 1
transform 1 0 47748 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_503
timestamp 1
transform 1 0 48300 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_505
timestamp 1636968456
transform 1 0 48484 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_517
timestamp 1636968456
transform 1 0 49588 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_529
timestamp 1636968456
transform 1 0 50692 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_541
timestamp 1636968456
transform 1 0 51796 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_553
timestamp 1
transform 1 0 52900 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_559
timestamp 1
transform 1 0 53452 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_561
timestamp 1636968456
transform 1 0 53636 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_573
timestamp 1636968456
transform 1 0 54740 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_585
timestamp 1636968456
transform 1 0 55844 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_597
timestamp 1636968456
transform 1 0 56948 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_609
timestamp 1
transform 1 0 58052 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_615
timestamp 1
transform 1 0 58604 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_617
timestamp 1636968456
transform 1 0 58788 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_629
timestamp 1636968456
transform 1 0 59892 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_641
timestamp 1636968456
transform 1 0 60996 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_653
timestamp 1636968456
transform 1 0 62100 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_665
timestamp 1
transform 1 0 63204 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_671
timestamp 1
transform 1 0 63756 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_673
timestamp 1636968456
transform 1 0 63940 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_685
timestamp 1636968456
transform 1 0 65044 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_697
timestamp 1636968456
transform 1 0 66148 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_709
timestamp 1636968456
transform 1 0 67252 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_721
timestamp 1
transform 1 0 68356 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_727
timestamp 1
transform 1 0 68908 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_729
timestamp 1636968456
transform 1 0 69092 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_741
timestamp 1636968456
transform 1 0 70196 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_753
timestamp 1636968456
transform 1 0 71300 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_765
timestamp 1636968456
transform 1 0 72404 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_777
timestamp 1
transform 1 0 73508 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_783
timestamp 1
transform 1 0 74060 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_785
timestamp 1636968456
transform 1 0 74244 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_797
timestamp 1636968456
transform 1 0 75348 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_809
timestamp 1636968456
transform 1 0 76452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_115_821
timestamp 1
transform 1 0 77556 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1636968456
transform 1 0 2300 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1636968456
transform 1 0 3404 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1
transform 1 0 4508 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1636968456
transform 1 0 4692 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_41
timestamp 1636968456
transform 1 0 5796 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_53
timestamp 1636968456
transform 1 0 6900 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_65
timestamp 1636968456
transform 1 0 8004 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_77
timestamp 1
transform 1 0 9108 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1
transform 1 0 9660 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_85
timestamp 1636968456
transform 1 0 9844 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_97
timestamp 1636968456
transform 1 0 10948 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_109
timestamp 1636968456
transform 1 0 12052 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_121
timestamp 1636968456
transform 1 0 13156 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_133
timestamp 1
transform 1 0 14260 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_139
timestamp 1
transform 1 0 14812 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_141
timestamp 1636968456
transform 1 0 14996 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_153
timestamp 1636968456
transform 1 0 16100 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_165
timestamp 1636968456
transform 1 0 17204 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_177
timestamp 1636968456
transform 1 0 18308 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_189
timestamp 1
transform 1 0 19412 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_195
timestamp 1
transform 1 0 19964 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_197
timestamp 1636968456
transform 1 0 20148 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_209
timestamp 1636968456
transform 1 0 21252 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_221
timestamp 1636968456
transform 1 0 22356 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_233
timestamp 1636968456
transform 1 0 23460 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_245
timestamp 1
transform 1 0 24564 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_251
timestamp 1
transform 1 0 25116 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_253
timestamp 1636968456
transform 1 0 25300 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_265
timestamp 1636968456
transform 1 0 26404 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_277
timestamp 1636968456
transform 1 0 27508 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_289
timestamp 1636968456
transform 1 0 28612 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_301
timestamp 1
transform 1 0 29716 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_307
timestamp 1
transform 1 0 30268 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_309
timestamp 1636968456
transform 1 0 30452 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_321
timestamp 1636968456
transform 1 0 31556 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_333
timestamp 1636968456
transform 1 0 32660 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_345
timestamp 1636968456
transform 1 0 33764 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_357
timestamp 1
transform 1 0 34868 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_363
timestamp 1
transform 1 0 35420 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_365
timestamp 1636968456
transform 1 0 35604 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_377
timestamp 1636968456
transform 1 0 36708 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_389
timestamp 1636968456
transform 1 0 37812 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_401
timestamp 1636968456
transform 1 0 38916 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_413
timestamp 1
transform 1 0 40020 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_419
timestamp 1
transform 1 0 40572 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_421
timestamp 1636968456
transform 1 0 40756 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_433
timestamp 1636968456
transform 1 0 41860 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_445
timestamp 1636968456
transform 1 0 42964 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_457
timestamp 1636968456
transform 1 0 44068 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_469
timestamp 1
transform 1 0 45172 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_475
timestamp 1
transform 1 0 45724 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_477
timestamp 1636968456
transform 1 0 45908 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_489
timestamp 1636968456
transform 1 0 47012 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_501
timestamp 1636968456
transform 1 0 48116 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_513
timestamp 1636968456
transform 1 0 49220 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_525
timestamp 1
transform 1 0 50324 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_531
timestamp 1
transform 1 0 50876 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_533
timestamp 1636968456
transform 1 0 51060 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_545
timestamp 1636968456
transform 1 0 52164 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_557
timestamp 1636968456
transform 1 0 53268 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_569
timestamp 1636968456
transform 1 0 54372 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_581
timestamp 1
transform 1 0 55476 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_587
timestamp 1
transform 1 0 56028 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_589
timestamp 1636968456
transform 1 0 56212 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_601
timestamp 1636968456
transform 1 0 57316 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_613
timestamp 1636968456
transform 1 0 58420 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_625
timestamp 1636968456
transform 1 0 59524 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_637
timestamp 1
transform 1 0 60628 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_643
timestamp 1
transform 1 0 61180 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_645
timestamp 1636968456
transform 1 0 61364 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_657
timestamp 1636968456
transform 1 0 62468 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_669
timestamp 1636968456
transform 1 0 63572 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_681
timestamp 1636968456
transform 1 0 64676 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_693
timestamp 1
transform 1 0 65780 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_699
timestamp 1
transform 1 0 66332 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_701
timestamp 1636968456
transform 1 0 66516 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_713
timestamp 1636968456
transform 1 0 67620 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_725
timestamp 1636968456
transform 1 0 68724 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_737
timestamp 1636968456
transform 1 0 69828 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_749
timestamp 1
transform 1 0 70932 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_755
timestamp 1
transform 1 0 71484 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_757
timestamp 1636968456
transform 1 0 71668 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_769
timestamp 1636968456
transform 1 0 72772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_781
timestamp 1636968456
transform 1 0 73876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_793
timestamp 1636968456
transform 1 0 74980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_805
timestamp 1
transform 1 0 76084 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_811
timestamp 1
transform 1 0 76636 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_813
timestamp 1
transform 1 0 76820 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_116_821
timestamp 1
transform 1 0 77556 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1636968456
transform 1 0 2300 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1636968456
transform 1 0 3404 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_27
timestamp 1636968456
transform 1 0 4508 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_39
timestamp 1636968456
transform 1 0 5612 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_51
timestamp 1
transform 1 0 6716 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_55
timestamp 1
transform 1 0 7084 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_57
timestamp 1636968456
transform 1 0 7268 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_69
timestamp 1636968456
transform 1 0 8372 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_81
timestamp 1636968456
transform 1 0 9476 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_93
timestamp 1636968456
transform 1 0 10580 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_105
timestamp 1
transform 1 0 11684 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_111
timestamp 1
transform 1 0 12236 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_113
timestamp 1636968456
transform 1 0 12420 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_125
timestamp 1636968456
transform 1 0 13524 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_137
timestamp 1636968456
transform 1 0 14628 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_149
timestamp 1636968456
transform 1 0 15732 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_161
timestamp 1
transform 1 0 16836 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_167
timestamp 1
transform 1 0 17388 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_169
timestamp 1636968456
transform 1 0 17572 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_181
timestamp 1636968456
transform 1 0 18676 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_193
timestamp 1636968456
transform 1 0 19780 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_205
timestamp 1636968456
transform 1 0 20884 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_217
timestamp 1
transform 1 0 21988 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_223
timestamp 1
transform 1 0 22540 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_225
timestamp 1636968456
transform 1 0 22724 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_237
timestamp 1636968456
transform 1 0 23828 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_249
timestamp 1636968456
transform 1 0 24932 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_261
timestamp 1636968456
transform 1 0 26036 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_273
timestamp 1
transform 1 0 27140 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_279
timestamp 1
transform 1 0 27692 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_281
timestamp 1636968456
transform 1 0 27876 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_293
timestamp 1636968456
transform 1 0 28980 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_305
timestamp 1636968456
transform 1 0 30084 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_317
timestamp 1636968456
transform 1 0 31188 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_329
timestamp 1
transform 1 0 32292 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_335
timestamp 1
transform 1 0 32844 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_337
timestamp 1636968456
transform 1 0 33028 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_349
timestamp 1636968456
transform 1 0 34132 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_361
timestamp 1636968456
transform 1 0 35236 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_373
timestamp 1636968456
transform 1 0 36340 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_385
timestamp 1
transform 1 0 37444 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_391
timestamp 1
transform 1 0 37996 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_393
timestamp 1636968456
transform 1 0 38180 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_405
timestamp 1636968456
transform 1 0 39284 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_417
timestamp 1636968456
transform 1 0 40388 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_429
timestamp 1636968456
transform 1 0 41492 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_441
timestamp 1
transform 1 0 42596 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_447
timestamp 1
transform 1 0 43148 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_449
timestamp 1636968456
transform 1 0 43332 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_461
timestamp 1636968456
transform 1 0 44436 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_473
timestamp 1636968456
transform 1 0 45540 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_485
timestamp 1636968456
transform 1 0 46644 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_497
timestamp 1
transform 1 0 47748 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_503
timestamp 1
transform 1 0 48300 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_505
timestamp 1636968456
transform 1 0 48484 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_517
timestamp 1636968456
transform 1 0 49588 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_529
timestamp 1636968456
transform 1 0 50692 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_541
timestamp 1636968456
transform 1 0 51796 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_553
timestamp 1
transform 1 0 52900 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_559
timestamp 1
transform 1 0 53452 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_561
timestamp 1636968456
transform 1 0 53636 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_573
timestamp 1636968456
transform 1 0 54740 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_585
timestamp 1636968456
transform 1 0 55844 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_597
timestamp 1636968456
transform 1 0 56948 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_609
timestamp 1
transform 1 0 58052 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_615
timestamp 1
transform 1 0 58604 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_617
timestamp 1636968456
transform 1 0 58788 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_629
timestamp 1636968456
transform 1 0 59892 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_641
timestamp 1636968456
transform 1 0 60996 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_653
timestamp 1636968456
transform 1 0 62100 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_665
timestamp 1
transform 1 0 63204 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_671
timestamp 1
transform 1 0 63756 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_673
timestamp 1636968456
transform 1 0 63940 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_685
timestamp 1636968456
transform 1 0 65044 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_697
timestamp 1636968456
transform 1 0 66148 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_709
timestamp 1636968456
transform 1 0 67252 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_721
timestamp 1
transform 1 0 68356 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_727
timestamp 1
transform 1 0 68908 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_729
timestamp 1636968456
transform 1 0 69092 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_741
timestamp 1636968456
transform 1 0 70196 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_753
timestamp 1636968456
transform 1 0 71300 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_765
timestamp 1636968456
transform 1 0 72404 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_777
timestamp 1
transform 1 0 73508 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_783
timestamp 1
transform 1 0 74060 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_785
timestamp 1636968456
transform 1 0 74244 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_797
timestamp 1636968456
transform 1 0 75348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_809
timestamp 1636968456
transform 1 0 76452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_117_821
timestamp 1
transform 1 0 77556 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1636968456
transform 1 0 2300 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1636968456
transform 1 0 3404 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1
transform 1 0 4508 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1636968456
transform 1 0 4692 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_41
timestamp 1636968456
transform 1 0 5796 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_53
timestamp 1636968456
transform 1 0 6900 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_65
timestamp 1636968456
transform 1 0 8004 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1
transform 1 0 9108 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1
transform 1 0 9660 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_85
timestamp 1636968456
transform 1 0 9844 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_97
timestamp 1636968456
transform 1 0 10948 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_109
timestamp 1636968456
transform 1 0 12052 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_121
timestamp 1636968456
transform 1 0 13156 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1
transform 1 0 14260 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1
transform 1 0 14812 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_141
timestamp 1636968456
transform 1 0 14996 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_153
timestamp 1636968456
transform 1 0 16100 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_165
timestamp 1636968456
transform 1 0 17204 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_177
timestamp 1636968456
transform 1 0 18308 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1
transform 1 0 19412 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1
transform 1 0 19964 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_197
timestamp 1636968456
transform 1 0 20148 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_209
timestamp 1636968456
transform 1 0 21252 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_221
timestamp 1636968456
transform 1 0 22356 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_233
timestamp 1636968456
transform 1 0 23460 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_245
timestamp 1
transform 1 0 24564 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1
transform 1 0 25116 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_253
timestamp 1636968456
transform 1 0 25300 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_265
timestamp 1636968456
transform 1 0 26404 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_277
timestamp 1636968456
transform 1 0 27508 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_289
timestamp 1636968456
transform 1 0 28612 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_301
timestamp 1
transform 1 0 29716 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_307
timestamp 1
transform 1 0 30268 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_309
timestamp 1636968456
transform 1 0 30452 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_321
timestamp 1636968456
transform 1 0 31556 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_333
timestamp 1636968456
transform 1 0 32660 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_345
timestamp 1636968456
transform 1 0 33764 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_357
timestamp 1
transform 1 0 34868 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_363
timestamp 1
transform 1 0 35420 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_365
timestamp 1636968456
transform 1 0 35604 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_377
timestamp 1636968456
transform 1 0 36708 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_389
timestamp 1636968456
transform 1 0 37812 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_401
timestamp 1636968456
transform 1 0 38916 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_413
timestamp 1
transform 1 0 40020 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1
transform 1 0 40572 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_421
timestamp 1636968456
transform 1 0 40756 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_433
timestamp 1636968456
transform 1 0 41860 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_445
timestamp 1636968456
transform 1 0 42964 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_457
timestamp 1636968456
transform 1 0 44068 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_469
timestamp 1
transform 1 0 45172 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_475
timestamp 1
transform 1 0 45724 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_477
timestamp 1636968456
transform 1 0 45908 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_489
timestamp 1636968456
transform 1 0 47012 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_501
timestamp 1636968456
transform 1 0 48116 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_513
timestamp 1636968456
transform 1 0 49220 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_525
timestamp 1
transform 1 0 50324 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_531
timestamp 1
transform 1 0 50876 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_533
timestamp 1636968456
transform 1 0 51060 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_545
timestamp 1636968456
transform 1 0 52164 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_557
timestamp 1636968456
transform 1 0 53268 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_569
timestamp 1636968456
transform 1 0 54372 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_581
timestamp 1
transform 1 0 55476 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1
transform 1 0 56028 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_589
timestamp 1636968456
transform 1 0 56212 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_601
timestamp 1636968456
transform 1 0 57316 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_613
timestamp 1636968456
transform 1 0 58420 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_625
timestamp 1636968456
transform 1 0 59524 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_637
timestamp 1
transform 1 0 60628 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_643
timestamp 1
transform 1 0 61180 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_645
timestamp 1636968456
transform 1 0 61364 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_657
timestamp 1636968456
transform 1 0 62468 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_669
timestamp 1636968456
transform 1 0 63572 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_681
timestamp 1636968456
transform 1 0 64676 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_693
timestamp 1
transform 1 0 65780 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1
transform 1 0 66332 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_701
timestamp 1636968456
transform 1 0 66516 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_713
timestamp 1636968456
transform 1 0 67620 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_725
timestamp 1636968456
transform 1 0 68724 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_737
timestamp 1636968456
transform 1 0 69828 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_749
timestamp 1
transform 1 0 70932 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_755
timestamp 1
transform 1 0 71484 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_757
timestamp 1636968456
transform 1 0 71668 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_769
timestamp 1636968456
transform 1 0 72772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_781
timestamp 1636968456
transform 1 0 73876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_793
timestamp 1636968456
transform 1 0 74980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_805
timestamp 1
transform 1 0 76084 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_811
timestamp 1
transform 1 0 76636 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_813
timestamp 1
transform 1 0 76820 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_821
timestamp 1
transform 1 0 77556 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1636968456
transform 1 0 2300 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1636968456
transform 1 0 3404 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_27
timestamp 1636968456
transform 1 0 4508 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_39
timestamp 1636968456
transform 1 0 5612 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1
transform 1 0 6716 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1
transform 1 0 7084 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_57
timestamp 1636968456
transform 1 0 7268 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_69
timestamp 1636968456
transform 1 0 8372 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_81
timestamp 1636968456
transform 1 0 9476 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_93
timestamp 1636968456
transform 1 0 10580 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1
transform 1 0 11684 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1
transform 1 0 12236 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_113
timestamp 1636968456
transform 1 0 12420 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_125
timestamp 1636968456
transform 1 0 13524 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_137
timestamp 1636968456
transform 1 0 14628 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_149
timestamp 1636968456
transform 1 0 15732 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1
transform 1 0 16836 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1
transform 1 0 17388 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_169
timestamp 1636968456
transform 1 0 17572 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_181
timestamp 1636968456
transform 1 0 18676 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_193
timestamp 1636968456
transform 1 0 19780 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_205
timestamp 1636968456
transform 1 0 20884 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_217
timestamp 1
transform 1 0 21988 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1
transform 1 0 22540 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_225
timestamp 1636968456
transform 1 0 22724 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_237
timestamp 1636968456
transform 1 0 23828 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_249
timestamp 1636968456
transform 1 0 24932 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_261
timestamp 1636968456
transform 1 0 26036 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_273
timestamp 1
transform 1 0 27140 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1
transform 1 0 27692 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_281
timestamp 1636968456
transform 1 0 27876 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_293
timestamp 1636968456
transform 1 0 28980 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_305
timestamp 1636968456
transform 1 0 30084 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_317
timestamp 1636968456
transform 1 0 31188 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_329
timestamp 1
transform 1 0 32292 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_335
timestamp 1
transform 1 0 32844 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_337
timestamp 1636968456
transform 1 0 33028 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_349
timestamp 1636968456
transform 1 0 34132 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_361
timestamp 1636968456
transform 1 0 35236 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_373
timestamp 1636968456
transform 1 0 36340 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_385
timestamp 1
transform 1 0 37444 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_391
timestamp 1
transform 1 0 37996 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_393
timestamp 1636968456
transform 1 0 38180 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_405
timestamp 1636968456
transform 1 0 39284 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_417
timestamp 1636968456
transform 1 0 40388 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_429
timestamp 1636968456
transform 1 0 41492 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_441
timestamp 1
transform 1 0 42596 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_447
timestamp 1
transform 1 0 43148 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_449
timestamp 1636968456
transform 1 0 43332 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_461
timestamp 1636968456
transform 1 0 44436 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_473
timestamp 1636968456
transform 1 0 45540 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_485
timestamp 1636968456
transform 1 0 46644 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_497
timestamp 1
transform 1 0 47748 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1
transform 1 0 48300 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_505
timestamp 1636968456
transform 1 0 48484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_517
timestamp 1636968456
transform 1 0 49588 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_529
timestamp 1636968456
transform 1 0 50692 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_541
timestamp 1636968456
transform 1 0 51796 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_553
timestamp 1
transform 1 0 52900 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_559
timestamp 1
transform 1 0 53452 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_561
timestamp 1636968456
transform 1 0 53636 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_573
timestamp 1636968456
transform 1 0 54740 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_585
timestamp 1636968456
transform 1 0 55844 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_597
timestamp 1636968456
transform 1 0 56948 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_609
timestamp 1
transform 1 0 58052 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_615
timestamp 1
transform 1 0 58604 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_617
timestamp 1636968456
transform 1 0 58788 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_629
timestamp 1636968456
transform 1 0 59892 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_641
timestamp 1636968456
transform 1 0 60996 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_653
timestamp 1636968456
transform 1 0 62100 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_665
timestamp 1
transform 1 0 63204 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_671
timestamp 1
transform 1 0 63756 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_673
timestamp 1636968456
transform 1 0 63940 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_685
timestamp 1636968456
transform 1 0 65044 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_697
timestamp 1636968456
transform 1 0 66148 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_709
timestamp 1636968456
transform 1 0 67252 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_721
timestamp 1
transform 1 0 68356 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_727
timestamp 1
transform 1 0 68908 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_729
timestamp 1636968456
transform 1 0 69092 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_741
timestamp 1636968456
transform 1 0 70196 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_753
timestamp 1636968456
transform 1 0 71300 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_765
timestamp 1636968456
transform 1 0 72404 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_777
timestamp 1
transform 1 0 73508 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_783
timestamp 1
transform 1 0 74060 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_785
timestamp 1636968456
transform 1 0 74244 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_797
timestamp 1636968456
transform 1 0 75348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_809
timestamp 1636968456
transform 1 0 76452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_119_821
timestamp 1
transform 1 0 77556 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_3
timestamp 1636968456
transform 1 0 2300 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_15
timestamp 1636968456
transform 1 0 3404 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1
transform 1 0 4508 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1636968456
transform 1 0 4692 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_41
timestamp 1636968456
transform 1 0 5796 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_53
timestamp 1636968456
transform 1 0 6900 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_65
timestamp 1636968456
transform 1 0 8004 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1
transform 1 0 9108 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1
transform 1 0 9660 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_85
timestamp 1636968456
transform 1 0 9844 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_97
timestamp 1636968456
transform 1 0 10948 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_109
timestamp 1636968456
transform 1 0 12052 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_121
timestamp 1636968456
transform 1 0 13156 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_133
timestamp 1
transform 1 0 14260 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1
transform 1 0 14812 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_141
timestamp 1636968456
transform 1 0 14996 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_153
timestamp 1636968456
transform 1 0 16100 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_165
timestamp 1636968456
transform 1 0 17204 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_177
timestamp 1636968456
transform 1 0 18308 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_189
timestamp 1
transform 1 0 19412 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_195
timestamp 1
transform 1 0 19964 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_197
timestamp 1636968456
transform 1 0 20148 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_209
timestamp 1636968456
transform 1 0 21252 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_221
timestamp 1636968456
transform 1 0 22356 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_233
timestamp 1636968456
transform 1 0 23460 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1
transform 1 0 24564 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1
transform 1 0 25116 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_253
timestamp 1636968456
transform 1 0 25300 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_265
timestamp 1636968456
transform 1 0 26404 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_277
timestamp 1636968456
transform 1 0 27508 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_289
timestamp 1636968456
transform 1 0 28612 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_301
timestamp 1
transform 1 0 29716 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_307
timestamp 1
transform 1 0 30268 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_309
timestamp 1636968456
transform 1 0 30452 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_321
timestamp 1636968456
transform 1 0 31556 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_333
timestamp 1636968456
transform 1 0 32660 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_345
timestamp 1636968456
transform 1 0 33764 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_357
timestamp 1
transform 1 0 34868 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1
transform 1 0 35420 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_365
timestamp 1636968456
transform 1 0 35604 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_377
timestamp 1636968456
transform 1 0 36708 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_389
timestamp 1636968456
transform 1 0 37812 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_401
timestamp 1636968456
transform 1 0 38916 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_413
timestamp 1
transform 1 0 40020 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_419
timestamp 1
transform 1 0 40572 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_421
timestamp 1636968456
transform 1 0 40756 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_433
timestamp 1636968456
transform 1 0 41860 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_445
timestamp 1636968456
transform 1 0 42964 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_457
timestamp 1636968456
transform 1 0 44068 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_469
timestamp 1
transform 1 0 45172 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_475
timestamp 1
transform 1 0 45724 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_477
timestamp 1636968456
transform 1 0 45908 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_489
timestamp 1636968456
transform 1 0 47012 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_501
timestamp 1636968456
transform 1 0 48116 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_513
timestamp 1636968456
transform 1 0 49220 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_525
timestamp 1
transform 1 0 50324 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_531
timestamp 1
transform 1 0 50876 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_533
timestamp 1636968456
transform 1 0 51060 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_545
timestamp 1636968456
transform 1 0 52164 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_557
timestamp 1636968456
transform 1 0 53268 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_569
timestamp 1636968456
transform 1 0 54372 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_581
timestamp 1
transform 1 0 55476 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_587
timestamp 1
transform 1 0 56028 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_589
timestamp 1636968456
transform 1 0 56212 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_601
timestamp 1636968456
transform 1 0 57316 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_613
timestamp 1636968456
transform 1 0 58420 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_625
timestamp 1636968456
transform 1 0 59524 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_637
timestamp 1
transform 1 0 60628 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_643
timestamp 1
transform 1 0 61180 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_645
timestamp 1636968456
transform 1 0 61364 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_657
timestamp 1636968456
transform 1 0 62468 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_669
timestamp 1636968456
transform 1 0 63572 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_681
timestamp 1636968456
transform 1 0 64676 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_693
timestamp 1
transform 1 0 65780 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_699
timestamp 1
transform 1 0 66332 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_701
timestamp 1636968456
transform 1 0 66516 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_713
timestamp 1636968456
transform 1 0 67620 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_725
timestamp 1636968456
transform 1 0 68724 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_737
timestamp 1636968456
transform 1 0 69828 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_749
timestamp 1
transform 1 0 70932 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_755
timestamp 1
transform 1 0 71484 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_757
timestamp 1636968456
transform 1 0 71668 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_769
timestamp 1636968456
transform 1 0 72772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_781
timestamp 1636968456
transform 1 0 73876 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_793
timestamp 1636968456
transform 1 0 74980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_805
timestamp 1
transform 1 0 76084 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_811
timestamp 1
transform 1 0 76636 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_813
timestamp 1
transform 1 0 76820 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_821
timestamp 1
transform 1 0 77556 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1636968456
transform 1 0 2300 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1636968456
transform 1 0 3404 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_27
timestamp 1636968456
transform 1 0 4508 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_39
timestamp 1636968456
transform 1 0 5612 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1
transform 1 0 6716 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1
transform 1 0 7084 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_57
timestamp 1636968456
transform 1 0 7268 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_69
timestamp 1636968456
transform 1 0 8372 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_81
timestamp 1636968456
transform 1 0 9476 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_93
timestamp 1636968456
transform 1 0 10580 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1
transform 1 0 11684 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1
transform 1 0 12236 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_113
timestamp 1636968456
transform 1 0 12420 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_125
timestamp 1636968456
transform 1 0 13524 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_137
timestamp 1636968456
transform 1 0 14628 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_149
timestamp 1636968456
transform 1 0 15732 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1
transform 1 0 16836 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1
transform 1 0 17388 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_169
timestamp 1636968456
transform 1 0 17572 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_181
timestamp 1636968456
transform 1 0 18676 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_193
timestamp 1636968456
transform 1 0 19780 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_205
timestamp 1636968456
transform 1 0 20884 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_217
timestamp 1
transform 1 0 21988 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_223
timestamp 1
transform 1 0 22540 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_225
timestamp 1636968456
transform 1 0 22724 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_237
timestamp 1636968456
transform 1 0 23828 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_249
timestamp 1636968456
transform 1 0 24932 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_261
timestamp 1636968456
transform 1 0 26036 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_273
timestamp 1
transform 1 0 27140 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1
transform 1 0 27692 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_281
timestamp 1636968456
transform 1 0 27876 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_293
timestamp 1636968456
transform 1 0 28980 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_305
timestamp 1636968456
transform 1 0 30084 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_317
timestamp 1636968456
transform 1 0 31188 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_329
timestamp 1
transform 1 0 32292 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_335
timestamp 1
transform 1 0 32844 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_337
timestamp 1636968456
transform 1 0 33028 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_349
timestamp 1636968456
transform 1 0 34132 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_361
timestamp 1636968456
transform 1 0 35236 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_373
timestamp 1636968456
transform 1 0 36340 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_385
timestamp 1
transform 1 0 37444 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_391
timestamp 1
transform 1 0 37996 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_393
timestamp 1636968456
transform 1 0 38180 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_405
timestamp 1636968456
transform 1 0 39284 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_417
timestamp 1636968456
transform 1 0 40388 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_429
timestamp 1636968456
transform 1 0 41492 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_441
timestamp 1
transform 1 0 42596 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_447
timestamp 1
transform 1 0 43148 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_449
timestamp 1636968456
transform 1 0 43332 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_461
timestamp 1636968456
transform 1 0 44436 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_473
timestamp 1636968456
transform 1 0 45540 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_485
timestamp 1636968456
transform 1 0 46644 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_497
timestamp 1
transform 1 0 47748 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_503
timestamp 1
transform 1 0 48300 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_505
timestamp 1636968456
transform 1 0 48484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_517
timestamp 1636968456
transform 1 0 49588 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_529
timestamp 1636968456
transform 1 0 50692 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_541
timestamp 1636968456
transform 1 0 51796 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_553
timestamp 1
transform 1 0 52900 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_559
timestamp 1
transform 1 0 53452 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_561
timestamp 1636968456
transform 1 0 53636 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_573
timestamp 1636968456
transform 1 0 54740 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_585
timestamp 1636968456
transform 1 0 55844 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_597
timestamp 1636968456
transform 1 0 56948 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_609
timestamp 1
transform 1 0 58052 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_615
timestamp 1
transform 1 0 58604 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_617
timestamp 1636968456
transform 1 0 58788 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_629
timestamp 1636968456
transform 1 0 59892 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_641
timestamp 1636968456
transform 1 0 60996 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_653
timestamp 1636968456
transform 1 0 62100 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_665
timestamp 1
transform 1 0 63204 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_671
timestamp 1
transform 1 0 63756 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_673
timestamp 1636968456
transform 1 0 63940 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_685
timestamp 1636968456
transform 1 0 65044 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_697
timestamp 1636968456
transform 1 0 66148 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_709
timestamp 1636968456
transform 1 0 67252 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_721
timestamp 1
transform 1 0 68356 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_727
timestamp 1
transform 1 0 68908 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_729
timestamp 1636968456
transform 1 0 69092 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_741
timestamp 1636968456
transform 1 0 70196 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_753
timestamp 1636968456
transform 1 0 71300 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_765
timestamp 1636968456
transform 1 0 72404 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_777
timestamp 1
transform 1 0 73508 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_783
timestamp 1
transform 1 0 74060 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_785
timestamp 1636968456
transform 1 0 74244 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_797
timestamp 1636968456
transform 1 0 75348 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_809
timestamp 1636968456
transform 1 0 76452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_121_821
timestamp 1
transform 1 0 77556 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_3
timestamp 1636968456
transform 1 0 2300 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_15
timestamp 1636968456
transform 1 0 3404 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1
transform 1 0 4508 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1636968456
transform 1 0 4692 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_41
timestamp 1636968456
transform 1 0 5796 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_53
timestamp 1636968456
transform 1 0 6900 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_65
timestamp 1636968456
transform 1 0 8004 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1
transform 1 0 9108 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1
transform 1 0 9660 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_85
timestamp 1636968456
transform 1 0 9844 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_97
timestamp 1636968456
transform 1 0 10948 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_109
timestamp 1636968456
transform 1 0 12052 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_121
timestamp 1636968456
transform 1 0 13156 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_133
timestamp 1
transform 1 0 14260 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_139
timestamp 1
transform 1 0 14812 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_141
timestamp 1636968456
transform 1 0 14996 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_153
timestamp 1636968456
transform 1 0 16100 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_165
timestamp 1636968456
transform 1 0 17204 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_177
timestamp 1636968456
transform 1 0 18308 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_189
timestamp 1
transform 1 0 19412 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_195
timestamp 1
transform 1 0 19964 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_197
timestamp 1636968456
transform 1 0 20148 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_209
timestamp 1636968456
transform 1 0 21252 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_221
timestamp 1636968456
transform 1 0 22356 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_233
timestamp 1636968456
transform 1 0 23460 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_245
timestamp 1
transform 1 0 24564 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_251
timestamp 1
transform 1 0 25116 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_253
timestamp 1636968456
transform 1 0 25300 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_265
timestamp 1636968456
transform 1 0 26404 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_277
timestamp 1636968456
transform 1 0 27508 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_289
timestamp 1636968456
transform 1 0 28612 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_301
timestamp 1
transform 1 0 29716 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_307
timestamp 1
transform 1 0 30268 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_309
timestamp 1636968456
transform 1 0 30452 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_321
timestamp 1636968456
transform 1 0 31556 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_333
timestamp 1636968456
transform 1 0 32660 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_345
timestamp 1636968456
transform 1 0 33764 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_357
timestamp 1
transform 1 0 34868 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_363
timestamp 1
transform 1 0 35420 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_365
timestamp 1636968456
transform 1 0 35604 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_377
timestamp 1636968456
transform 1 0 36708 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_389
timestamp 1636968456
transform 1 0 37812 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_401
timestamp 1636968456
transform 1 0 38916 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_413
timestamp 1
transform 1 0 40020 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_419
timestamp 1
transform 1 0 40572 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_421
timestamp 1636968456
transform 1 0 40756 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_433
timestamp 1636968456
transform 1 0 41860 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_445
timestamp 1636968456
transform 1 0 42964 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_457
timestamp 1636968456
transform 1 0 44068 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_469
timestamp 1
transform 1 0 45172 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_475
timestamp 1
transform 1 0 45724 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_477
timestamp 1636968456
transform 1 0 45908 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_489
timestamp 1636968456
transform 1 0 47012 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_501
timestamp 1636968456
transform 1 0 48116 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_513
timestamp 1636968456
transform 1 0 49220 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_525
timestamp 1
transform 1 0 50324 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_531
timestamp 1
transform 1 0 50876 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_533
timestamp 1636968456
transform 1 0 51060 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_545
timestamp 1636968456
transform 1 0 52164 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_557
timestamp 1636968456
transform 1 0 53268 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_569
timestamp 1636968456
transform 1 0 54372 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_581
timestamp 1
transform 1 0 55476 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_587
timestamp 1
transform 1 0 56028 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_589
timestamp 1636968456
transform 1 0 56212 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_601
timestamp 1636968456
transform 1 0 57316 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_613
timestamp 1636968456
transform 1 0 58420 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_625
timestamp 1636968456
transform 1 0 59524 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_637
timestamp 1
transform 1 0 60628 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_643
timestamp 1
transform 1 0 61180 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_645
timestamp 1636968456
transform 1 0 61364 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_657
timestamp 1636968456
transform 1 0 62468 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_669
timestamp 1636968456
transform 1 0 63572 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_681
timestamp 1636968456
transform 1 0 64676 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_693
timestamp 1
transform 1 0 65780 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_699
timestamp 1
transform 1 0 66332 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_701
timestamp 1636968456
transform 1 0 66516 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_713
timestamp 1636968456
transform 1 0 67620 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_725
timestamp 1636968456
transform 1 0 68724 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_737
timestamp 1636968456
transform 1 0 69828 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_749
timestamp 1
transform 1 0 70932 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_755
timestamp 1
transform 1 0 71484 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_757
timestamp 1636968456
transform 1 0 71668 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_769
timestamp 1636968456
transform 1 0 72772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_781
timestamp 1636968456
transform 1 0 73876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_793
timestamp 1636968456
transform 1 0 74980 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_805
timestamp 1
transform 1 0 76084 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_811
timestamp 1
transform 1 0 76636 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_813
timestamp 1
transform 1 0 76820 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_821
timestamp 1
transform 1 0 77556 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636968456
transform 1 0 2300 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636968456
transform 1 0 3404 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_27
timestamp 1636968456
transform 1 0 4508 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_39
timestamp 1636968456
transform 1 0 5612 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_51
timestamp 1
transform 1 0 6716 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1
transform 1 0 7084 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_57
timestamp 1636968456
transform 1 0 7268 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_69
timestamp 1636968456
transform 1 0 8372 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_81
timestamp 1636968456
transform 1 0 9476 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_93
timestamp 1636968456
transform 1 0 10580 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_105
timestamp 1
transform 1 0 11684 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_111
timestamp 1
transform 1 0 12236 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_113
timestamp 1636968456
transform 1 0 12420 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_125
timestamp 1636968456
transform 1 0 13524 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_137
timestamp 1636968456
transform 1 0 14628 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_149
timestamp 1636968456
transform 1 0 15732 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_161
timestamp 1
transform 1 0 16836 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_167
timestamp 1
transform 1 0 17388 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_169
timestamp 1636968456
transform 1 0 17572 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_181
timestamp 1636968456
transform 1 0 18676 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_193
timestamp 1636968456
transform 1 0 19780 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_205
timestamp 1636968456
transform 1 0 20884 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_217
timestamp 1
transform 1 0 21988 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_223
timestamp 1
transform 1 0 22540 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_225
timestamp 1636968456
transform 1 0 22724 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_237
timestamp 1636968456
transform 1 0 23828 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_249
timestamp 1636968456
transform 1 0 24932 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_261
timestamp 1636968456
transform 1 0 26036 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_273
timestamp 1
transform 1 0 27140 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_279
timestamp 1
transform 1 0 27692 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_281
timestamp 1636968456
transform 1 0 27876 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_293
timestamp 1636968456
transform 1 0 28980 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_305
timestamp 1636968456
transform 1 0 30084 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_317
timestamp 1636968456
transform 1 0 31188 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_329
timestamp 1
transform 1 0 32292 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_335
timestamp 1
transform 1 0 32844 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_337
timestamp 1636968456
transform 1 0 33028 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_349
timestamp 1636968456
transform 1 0 34132 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_361
timestamp 1636968456
transform 1 0 35236 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_373
timestamp 1636968456
transform 1 0 36340 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_385
timestamp 1
transform 1 0 37444 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_391
timestamp 1
transform 1 0 37996 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_393
timestamp 1636968456
transform 1 0 38180 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_405
timestamp 1636968456
transform 1 0 39284 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_417
timestamp 1636968456
transform 1 0 40388 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_429
timestamp 1636968456
transform 1 0 41492 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_441
timestamp 1
transform 1 0 42596 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_447
timestamp 1
transform 1 0 43148 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_449
timestamp 1636968456
transform 1 0 43332 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_461
timestamp 1636968456
transform 1 0 44436 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_473
timestamp 1636968456
transform 1 0 45540 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_485
timestamp 1636968456
transform 1 0 46644 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_497
timestamp 1
transform 1 0 47748 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_503
timestamp 1
transform 1 0 48300 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_505
timestamp 1636968456
transform 1 0 48484 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_517
timestamp 1636968456
transform 1 0 49588 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_529
timestamp 1636968456
transform 1 0 50692 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_541
timestamp 1636968456
transform 1 0 51796 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_553
timestamp 1
transform 1 0 52900 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_559
timestamp 1
transform 1 0 53452 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_561
timestamp 1636968456
transform 1 0 53636 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_573
timestamp 1636968456
transform 1 0 54740 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_585
timestamp 1636968456
transform 1 0 55844 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_597
timestamp 1636968456
transform 1 0 56948 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_609
timestamp 1
transform 1 0 58052 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_615
timestamp 1
transform 1 0 58604 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_617
timestamp 1636968456
transform 1 0 58788 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_629
timestamp 1636968456
transform 1 0 59892 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_641
timestamp 1636968456
transform 1 0 60996 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_653
timestamp 1636968456
transform 1 0 62100 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_665
timestamp 1
transform 1 0 63204 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_671
timestamp 1
transform 1 0 63756 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_673
timestamp 1636968456
transform 1 0 63940 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_685
timestamp 1636968456
transform 1 0 65044 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_697
timestamp 1636968456
transform 1 0 66148 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_709
timestamp 1636968456
transform 1 0 67252 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_721
timestamp 1
transform 1 0 68356 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_727
timestamp 1
transform 1 0 68908 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_729
timestamp 1636968456
transform 1 0 69092 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_741
timestamp 1636968456
transform 1 0 70196 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_753
timestamp 1636968456
transform 1 0 71300 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_765
timestamp 1636968456
transform 1 0 72404 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_777
timestamp 1
transform 1 0 73508 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_783
timestamp 1
transform 1 0 74060 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_785
timestamp 1636968456
transform 1 0 74244 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_797
timestamp 1636968456
transform 1 0 75348 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_809
timestamp 1636968456
transform 1 0 76452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_123_821
timestamp 1
transform 1 0 77556 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_3
timestamp 1636968456
transform 1 0 2300 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_15
timestamp 1636968456
transform 1 0 3404 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 1
transform 1 0 4508 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_29
timestamp 1636968456
transform 1 0 4692 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_41
timestamp 1636968456
transform 1 0 5796 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_53
timestamp 1636968456
transform 1 0 6900 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_65
timestamp 1636968456
transform 1 0 8004 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1
transform 1 0 9108 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1
transform 1 0 9660 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_85
timestamp 1636968456
transform 1 0 9844 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_97
timestamp 1636968456
transform 1 0 10948 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_109
timestamp 1636968456
transform 1 0 12052 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_121
timestamp 1636968456
transform 1 0 13156 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_133
timestamp 1
transform 1 0 14260 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_139
timestamp 1
transform 1 0 14812 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_141
timestamp 1636968456
transform 1 0 14996 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_153
timestamp 1636968456
transform 1 0 16100 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_165
timestamp 1636968456
transform 1 0 17204 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_177
timestamp 1636968456
transform 1 0 18308 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_189
timestamp 1
transform 1 0 19412 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_195
timestamp 1
transform 1 0 19964 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_197
timestamp 1636968456
transform 1 0 20148 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_209
timestamp 1636968456
transform 1 0 21252 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_221
timestamp 1636968456
transform 1 0 22356 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_233
timestamp 1636968456
transform 1 0 23460 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_245
timestamp 1
transform 1 0 24564 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_251
timestamp 1
transform 1 0 25116 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_253
timestamp 1636968456
transform 1 0 25300 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_265
timestamp 1636968456
transform 1 0 26404 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_277
timestamp 1636968456
transform 1 0 27508 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_289
timestamp 1636968456
transform 1 0 28612 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_301
timestamp 1
transform 1 0 29716 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_307
timestamp 1
transform 1 0 30268 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_309
timestamp 1636968456
transform 1 0 30452 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_321
timestamp 1636968456
transform 1 0 31556 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_333
timestamp 1636968456
transform 1 0 32660 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_345
timestamp 1636968456
transform 1 0 33764 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_357
timestamp 1
transform 1 0 34868 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_363
timestamp 1
transform 1 0 35420 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_365
timestamp 1636968456
transform 1 0 35604 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_377
timestamp 1636968456
transform 1 0 36708 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_389
timestamp 1636968456
transform 1 0 37812 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_401
timestamp 1636968456
transform 1 0 38916 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_413
timestamp 1
transform 1 0 40020 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_419
timestamp 1
transform 1 0 40572 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_421
timestamp 1636968456
transform 1 0 40756 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_433
timestamp 1636968456
transform 1 0 41860 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_445
timestamp 1636968456
transform 1 0 42964 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_457
timestamp 1636968456
transform 1 0 44068 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_469
timestamp 1
transform 1 0 45172 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_475
timestamp 1
transform 1 0 45724 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_477
timestamp 1636968456
transform 1 0 45908 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_489
timestamp 1636968456
transform 1 0 47012 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_501
timestamp 1636968456
transform 1 0 48116 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_513
timestamp 1636968456
transform 1 0 49220 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_525
timestamp 1
transform 1 0 50324 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_531
timestamp 1
transform 1 0 50876 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_533
timestamp 1636968456
transform 1 0 51060 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_545
timestamp 1636968456
transform 1 0 52164 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_557
timestamp 1636968456
transform 1 0 53268 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_569
timestamp 1636968456
transform 1 0 54372 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_581
timestamp 1
transform 1 0 55476 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_587
timestamp 1
transform 1 0 56028 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_589
timestamp 1636968456
transform 1 0 56212 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_601
timestamp 1636968456
transform 1 0 57316 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_613
timestamp 1636968456
transform 1 0 58420 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_625
timestamp 1636968456
transform 1 0 59524 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_637
timestamp 1
transform 1 0 60628 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_643
timestamp 1
transform 1 0 61180 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_645
timestamp 1636968456
transform 1 0 61364 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_657
timestamp 1636968456
transform 1 0 62468 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_669
timestamp 1636968456
transform 1 0 63572 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_681
timestamp 1636968456
transform 1 0 64676 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_693
timestamp 1
transform 1 0 65780 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_699
timestamp 1
transform 1 0 66332 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_701
timestamp 1636968456
transform 1 0 66516 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_713
timestamp 1636968456
transform 1 0 67620 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_725
timestamp 1636968456
transform 1 0 68724 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_737
timestamp 1636968456
transform 1 0 69828 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_749
timestamp 1
transform 1 0 70932 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_755
timestamp 1
transform 1 0 71484 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_757
timestamp 1636968456
transform 1 0 71668 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_769
timestamp 1636968456
transform 1 0 72772 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_781
timestamp 1636968456
transform 1 0 73876 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_793
timestamp 1636968456
transform 1 0 74980 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_805
timestamp 1
transform 1 0 76084 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_811
timestamp 1
transform 1 0 76636 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_813
timestamp 1
transform 1 0 76820 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_124_821
timestamp 1
transform 1 0 77556 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_3
timestamp 1636968456
transform 1 0 2300 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_15
timestamp 1636968456
transform 1 0 3404 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_27
timestamp 1636968456
transform 1 0 4508 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_39
timestamp 1636968456
transform 1 0 5612 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_51
timestamp 1
transform 1 0 6716 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1
transform 1 0 7084 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_57
timestamp 1636968456
transform 1 0 7268 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_69
timestamp 1636968456
transform 1 0 8372 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_81
timestamp 1636968456
transform 1 0 9476 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_93
timestamp 1636968456
transform 1 0 10580 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_105
timestamp 1
transform 1 0 11684 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_111
timestamp 1
transform 1 0 12236 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_113
timestamp 1636968456
transform 1 0 12420 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_125
timestamp 1636968456
transform 1 0 13524 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_137
timestamp 1636968456
transform 1 0 14628 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_149
timestamp 1636968456
transform 1 0 15732 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_161
timestamp 1
transform 1 0 16836 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_167
timestamp 1
transform 1 0 17388 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_169
timestamp 1636968456
transform 1 0 17572 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_181
timestamp 1636968456
transform 1 0 18676 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_193
timestamp 1636968456
transform 1 0 19780 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_205
timestamp 1636968456
transform 1 0 20884 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_217
timestamp 1
transform 1 0 21988 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_223
timestamp 1
transform 1 0 22540 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_225
timestamp 1636968456
transform 1 0 22724 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_237
timestamp 1636968456
transform 1 0 23828 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_249
timestamp 1636968456
transform 1 0 24932 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_261
timestamp 1636968456
transform 1 0 26036 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_273
timestamp 1
transform 1 0 27140 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_279
timestamp 1
transform 1 0 27692 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_281
timestamp 1636968456
transform 1 0 27876 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_293
timestamp 1636968456
transform 1 0 28980 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_305
timestamp 1636968456
transform 1 0 30084 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_317
timestamp 1636968456
transform 1 0 31188 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_329
timestamp 1
transform 1 0 32292 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_335
timestamp 1
transform 1 0 32844 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_337
timestamp 1636968456
transform 1 0 33028 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_349
timestamp 1636968456
transform 1 0 34132 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_361
timestamp 1636968456
transform 1 0 35236 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_373
timestamp 1636968456
transform 1 0 36340 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_385
timestamp 1
transform 1 0 37444 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_391
timestamp 1
transform 1 0 37996 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_393
timestamp 1636968456
transform 1 0 38180 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_405
timestamp 1636968456
transform 1 0 39284 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_417
timestamp 1636968456
transform 1 0 40388 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_429
timestamp 1636968456
transform 1 0 41492 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_441
timestamp 1
transform 1 0 42596 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_447
timestamp 1
transform 1 0 43148 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_449
timestamp 1636968456
transform 1 0 43332 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_461
timestamp 1636968456
transform 1 0 44436 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_473
timestamp 1636968456
transform 1 0 45540 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_485
timestamp 1636968456
transform 1 0 46644 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_497
timestamp 1
transform 1 0 47748 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_503
timestamp 1
transform 1 0 48300 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_505
timestamp 1636968456
transform 1 0 48484 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_517
timestamp 1636968456
transform 1 0 49588 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_529
timestamp 1636968456
transform 1 0 50692 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_541
timestamp 1636968456
transform 1 0 51796 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_553
timestamp 1
transform 1 0 52900 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_559
timestamp 1
transform 1 0 53452 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_561
timestamp 1636968456
transform 1 0 53636 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_573
timestamp 1636968456
transform 1 0 54740 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_585
timestamp 1636968456
transform 1 0 55844 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_597
timestamp 1636968456
transform 1 0 56948 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_609
timestamp 1
transform 1 0 58052 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_615
timestamp 1
transform 1 0 58604 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_617
timestamp 1636968456
transform 1 0 58788 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_629
timestamp 1636968456
transform 1 0 59892 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_641
timestamp 1636968456
transform 1 0 60996 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_653
timestamp 1636968456
transform 1 0 62100 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_665
timestamp 1
transform 1 0 63204 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_671
timestamp 1
transform 1 0 63756 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_673
timestamp 1636968456
transform 1 0 63940 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_685
timestamp 1636968456
transform 1 0 65044 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_697
timestamp 1636968456
transform 1 0 66148 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_709
timestamp 1636968456
transform 1 0 67252 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_721
timestamp 1
transform 1 0 68356 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_727
timestamp 1
transform 1 0 68908 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_729
timestamp 1636968456
transform 1 0 69092 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_741
timestamp 1636968456
transform 1 0 70196 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_753
timestamp 1636968456
transform 1 0 71300 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_765
timestamp 1636968456
transform 1 0 72404 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_777
timestamp 1
transform 1 0 73508 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_783
timestamp 1
transform 1 0 74060 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_785
timestamp 1636968456
transform 1 0 74244 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_797
timestamp 1636968456
transform 1 0 75348 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_809
timestamp 1636968456
transform 1 0 76452 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_821
timestamp 1
transform 1 0 77556 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1636968456
transform 1 0 2300 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1636968456
transform 1 0 3404 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 1
transform 1 0 4508 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1636968456
transform 1 0 4692 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_41
timestamp 1636968456
transform 1 0 5796 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_53
timestamp 1636968456
transform 1 0 6900 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_65
timestamp 1636968456
transform 1 0 8004 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1
transform 1 0 9108 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1
transform 1 0 9660 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_85
timestamp 1636968456
transform 1 0 9844 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_97
timestamp 1636968456
transform 1 0 10948 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_109
timestamp 1636968456
transform 1 0 12052 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_121
timestamp 1636968456
transform 1 0 13156 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_133
timestamp 1
transform 1 0 14260 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_139
timestamp 1
transform 1 0 14812 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_141
timestamp 1636968456
transform 1 0 14996 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_153
timestamp 1636968456
transform 1 0 16100 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_165
timestamp 1636968456
transform 1 0 17204 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_177
timestamp 1636968456
transform 1 0 18308 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_189
timestamp 1
transform 1 0 19412 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_195
timestamp 1
transform 1 0 19964 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_197
timestamp 1636968456
transform 1 0 20148 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_209
timestamp 1636968456
transform 1 0 21252 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_221
timestamp 1636968456
transform 1 0 22356 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_233
timestamp 1636968456
transform 1 0 23460 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_245
timestamp 1
transform 1 0 24564 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_251
timestamp 1
transform 1 0 25116 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_253
timestamp 1636968456
transform 1 0 25300 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_265
timestamp 1636968456
transform 1 0 26404 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_277
timestamp 1636968456
transform 1 0 27508 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_289
timestamp 1636968456
transform 1 0 28612 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_301
timestamp 1
transform 1 0 29716 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_307
timestamp 1
transform 1 0 30268 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_309
timestamp 1636968456
transform 1 0 30452 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_321
timestamp 1636968456
transform 1 0 31556 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_333
timestamp 1636968456
transform 1 0 32660 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_345
timestamp 1636968456
transform 1 0 33764 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_357
timestamp 1
transform 1 0 34868 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_363
timestamp 1
transform 1 0 35420 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_365
timestamp 1636968456
transform 1 0 35604 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_377
timestamp 1636968456
transform 1 0 36708 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_389
timestamp 1636968456
transform 1 0 37812 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_401
timestamp 1636968456
transform 1 0 38916 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_413
timestamp 1
transform 1 0 40020 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_419
timestamp 1
transform 1 0 40572 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_421
timestamp 1636968456
transform 1 0 40756 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_433
timestamp 1636968456
transform 1 0 41860 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_445
timestamp 1636968456
transform 1 0 42964 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_457
timestamp 1636968456
transform 1 0 44068 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_469
timestamp 1
transform 1 0 45172 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_475
timestamp 1
transform 1 0 45724 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_477
timestamp 1636968456
transform 1 0 45908 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_489
timestamp 1636968456
transform 1 0 47012 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_501
timestamp 1636968456
transform 1 0 48116 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_513
timestamp 1636968456
transform 1 0 49220 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_525
timestamp 1
transform 1 0 50324 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_531
timestamp 1
transform 1 0 50876 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_533
timestamp 1636968456
transform 1 0 51060 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_545
timestamp 1636968456
transform 1 0 52164 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_557
timestamp 1636968456
transform 1 0 53268 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_569
timestamp 1636968456
transform 1 0 54372 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_581
timestamp 1
transform 1 0 55476 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_587
timestamp 1
transform 1 0 56028 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_589
timestamp 1636968456
transform 1 0 56212 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_601
timestamp 1636968456
transform 1 0 57316 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_613
timestamp 1636968456
transform 1 0 58420 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_625
timestamp 1636968456
transform 1 0 59524 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_637
timestamp 1
transform 1 0 60628 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_643
timestamp 1
transform 1 0 61180 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_645
timestamp 1636968456
transform 1 0 61364 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_657
timestamp 1636968456
transform 1 0 62468 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_669
timestamp 1636968456
transform 1 0 63572 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_681
timestamp 1636968456
transform 1 0 64676 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_693
timestamp 1
transform 1 0 65780 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_699
timestamp 1
transform 1 0 66332 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_701
timestamp 1636968456
transform 1 0 66516 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_713
timestamp 1636968456
transform 1 0 67620 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_725
timestamp 1636968456
transform 1 0 68724 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_737
timestamp 1636968456
transform 1 0 69828 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_749
timestamp 1
transform 1 0 70932 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_755
timestamp 1
transform 1 0 71484 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_757
timestamp 1636968456
transform 1 0 71668 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_769
timestamp 1636968456
transform 1 0 72772 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_781
timestamp 1636968456
transform 1 0 73876 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_793
timestamp 1636968456
transform 1 0 74980 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_805
timestamp 1
transform 1 0 76084 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_811
timestamp 1
transform 1 0 76636 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_126_813
timestamp 1
transform 1 0 76820 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_126_821
timestamp 1
transform 1 0 77556 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_3
timestamp 1636968456
transform 1 0 2300 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_15
timestamp 1636968456
transform 1 0 3404 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_27
timestamp 1636968456
transform 1 0 4508 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_39
timestamp 1636968456
transform 1 0 5612 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_51
timestamp 1
transform 1 0 6716 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1
transform 1 0 7084 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_57
timestamp 1636968456
transform 1 0 7268 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_69
timestamp 1636968456
transform 1 0 8372 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_81
timestamp 1636968456
transform 1 0 9476 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_93
timestamp 1636968456
transform 1 0 10580 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_105
timestamp 1
transform 1 0 11684 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_111
timestamp 1
transform 1 0 12236 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_113
timestamp 1636968456
transform 1 0 12420 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_125
timestamp 1636968456
transform 1 0 13524 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_137
timestamp 1636968456
transform 1 0 14628 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_149
timestamp 1636968456
transform 1 0 15732 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_161
timestamp 1
transform 1 0 16836 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_167
timestamp 1
transform 1 0 17388 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_169
timestamp 1636968456
transform 1 0 17572 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_181
timestamp 1636968456
transform 1 0 18676 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_193
timestamp 1636968456
transform 1 0 19780 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_205
timestamp 1636968456
transform 1 0 20884 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_217
timestamp 1
transform 1 0 21988 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_223
timestamp 1
transform 1 0 22540 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_225
timestamp 1636968456
transform 1 0 22724 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_237
timestamp 1636968456
transform 1 0 23828 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_249
timestamp 1636968456
transform 1 0 24932 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_261
timestamp 1636968456
transform 1 0 26036 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_273
timestamp 1
transform 1 0 27140 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_279
timestamp 1
transform 1 0 27692 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_281
timestamp 1636968456
transform 1 0 27876 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_293
timestamp 1636968456
transform 1 0 28980 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_305
timestamp 1636968456
transform 1 0 30084 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_317
timestamp 1636968456
transform 1 0 31188 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_329
timestamp 1
transform 1 0 32292 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_335
timestamp 1
transform 1 0 32844 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_337
timestamp 1636968456
transform 1 0 33028 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_349
timestamp 1636968456
transform 1 0 34132 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_361
timestamp 1636968456
transform 1 0 35236 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_373
timestamp 1636968456
transform 1 0 36340 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_385
timestamp 1
transform 1 0 37444 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_391
timestamp 1
transform 1 0 37996 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_393
timestamp 1636968456
transform 1 0 38180 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_405
timestamp 1636968456
transform 1 0 39284 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_417
timestamp 1636968456
transform 1 0 40388 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_429
timestamp 1636968456
transform 1 0 41492 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_441
timestamp 1
transform 1 0 42596 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_447
timestamp 1
transform 1 0 43148 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_449
timestamp 1636968456
transform 1 0 43332 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_461
timestamp 1636968456
transform 1 0 44436 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_473
timestamp 1636968456
transform 1 0 45540 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_485
timestamp 1636968456
transform 1 0 46644 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_497
timestamp 1
transform 1 0 47748 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_503
timestamp 1
transform 1 0 48300 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_505
timestamp 1636968456
transform 1 0 48484 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_517
timestamp 1636968456
transform 1 0 49588 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_529
timestamp 1636968456
transform 1 0 50692 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_541
timestamp 1636968456
transform 1 0 51796 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_553
timestamp 1
transform 1 0 52900 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_559
timestamp 1
transform 1 0 53452 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_561
timestamp 1636968456
transform 1 0 53636 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_573
timestamp 1636968456
transform 1 0 54740 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_585
timestamp 1636968456
transform 1 0 55844 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_597
timestamp 1636968456
transform 1 0 56948 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_609
timestamp 1
transform 1 0 58052 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_615
timestamp 1
transform 1 0 58604 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_617
timestamp 1636968456
transform 1 0 58788 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_629
timestamp 1636968456
transform 1 0 59892 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_641
timestamp 1636968456
transform 1 0 60996 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_653
timestamp 1636968456
transform 1 0 62100 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_665
timestamp 1
transform 1 0 63204 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_671
timestamp 1
transform 1 0 63756 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_673
timestamp 1636968456
transform 1 0 63940 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_685
timestamp 1636968456
transform 1 0 65044 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_697
timestamp 1636968456
transform 1 0 66148 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_709
timestamp 1636968456
transform 1 0 67252 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_721
timestamp 1
transform 1 0 68356 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_727
timestamp 1
transform 1 0 68908 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_729
timestamp 1636968456
transform 1 0 69092 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_741
timestamp 1636968456
transform 1 0 70196 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_753
timestamp 1636968456
transform 1 0 71300 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_765
timestamp 1636968456
transform 1 0 72404 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_777
timestamp 1
transform 1 0 73508 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_783
timestamp 1
transform 1 0 74060 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_785
timestamp 1636968456
transform 1 0 74244 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_797
timestamp 1636968456
transform 1 0 75348 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_809
timestamp 1636968456
transform 1 0 76452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_127_821
timestamp 1
transform 1 0 77556 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_3
timestamp 1636968456
transform 1 0 2300 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_15
timestamp 1636968456
transform 1 0 3404 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 1
transform 1 0 4508 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_29
timestamp 1636968456
transform 1 0 4692 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_41
timestamp 1636968456
transform 1 0 5796 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_53
timestamp 1636968456
transform 1 0 6900 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_65
timestamp 1636968456
transform 1 0 8004 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1
transform 1 0 9108 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1
transform 1 0 9660 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_85
timestamp 1636968456
transform 1 0 9844 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_97
timestamp 1636968456
transform 1 0 10948 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_109
timestamp 1636968456
transform 1 0 12052 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_121
timestamp 1636968456
transform 1 0 13156 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_133
timestamp 1
transform 1 0 14260 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_139
timestamp 1
transform 1 0 14812 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_141
timestamp 1636968456
transform 1 0 14996 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_153
timestamp 1636968456
transform 1 0 16100 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_165
timestamp 1636968456
transform 1 0 17204 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_177
timestamp 1636968456
transform 1 0 18308 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_189
timestamp 1
transform 1 0 19412 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_195
timestamp 1
transform 1 0 19964 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_197
timestamp 1636968456
transform 1 0 20148 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_209
timestamp 1636968456
transform 1 0 21252 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_221
timestamp 1636968456
transform 1 0 22356 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_233
timestamp 1636968456
transform 1 0 23460 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_245
timestamp 1
transform 1 0 24564 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_251
timestamp 1
transform 1 0 25116 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_253
timestamp 1636968456
transform 1 0 25300 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_265
timestamp 1636968456
transform 1 0 26404 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_277
timestamp 1636968456
transform 1 0 27508 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_289
timestamp 1636968456
transform 1 0 28612 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_301
timestamp 1
transform 1 0 29716 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_307
timestamp 1
transform 1 0 30268 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_309
timestamp 1636968456
transform 1 0 30452 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_321
timestamp 1636968456
transform 1 0 31556 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_333
timestamp 1636968456
transform 1 0 32660 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_345
timestamp 1636968456
transform 1 0 33764 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_357
timestamp 1
transform 1 0 34868 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_363
timestamp 1
transform 1 0 35420 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_365
timestamp 1636968456
transform 1 0 35604 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_377
timestamp 1636968456
transform 1 0 36708 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_389
timestamp 1636968456
transform 1 0 37812 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_401
timestamp 1636968456
transform 1 0 38916 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_413
timestamp 1
transform 1 0 40020 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_419
timestamp 1
transform 1 0 40572 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_421
timestamp 1636968456
transform 1 0 40756 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_433
timestamp 1636968456
transform 1 0 41860 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_445
timestamp 1636968456
transform 1 0 42964 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_457
timestamp 1636968456
transform 1 0 44068 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_469
timestamp 1
transform 1 0 45172 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_475
timestamp 1
transform 1 0 45724 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_477
timestamp 1636968456
transform 1 0 45908 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_489
timestamp 1636968456
transform 1 0 47012 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_501
timestamp 1636968456
transform 1 0 48116 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_513
timestamp 1636968456
transform 1 0 49220 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_525
timestamp 1
transform 1 0 50324 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_531
timestamp 1
transform 1 0 50876 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_533
timestamp 1636968456
transform 1 0 51060 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_545
timestamp 1636968456
transform 1 0 52164 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_557
timestamp 1636968456
transform 1 0 53268 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_569
timestamp 1636968456
transform 1 0 54372 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_581
timestamp 1
transform 1 0 55476 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_587
timestamp 1
transform 1 0 56028 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_589
timestamp 1636968456
transform 1 0 56212 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_601
timestamp 1636968456
transform 1 0 57316 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_613
timestamp 1636968456
transform 1 0 58420 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_625
timestamp 1636968456
transform 1 0 59524 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_637
timestamp 1
transform 1 0 60628 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_643
timestamp 1
transform 1 0 61180 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_645
timestamp 1636968456
transform 1 0 61364 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_657
timestamp 1636968456
transform 1 0 62468 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_669
timestamp 1636968456
transform 1 0 63572 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_681
timestamp 1636968456
transform 1 0 64676 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_693
timestamp 1
transform 1 0 65780 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_699
timestamp 1
transform 1 0 66332 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_701
timestamp 1636968456
transform 1 0 66516 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_713
timestamp 1636968456
transform 1 0 67620 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_725
timestamp 1636968456
transform 1 0 68724 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_737
timestamp 1636968456
transform 1 0 69828 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_749
timestamp 1
transform 1 0 70932 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_755
timestamp 1
transform 1 0 71484 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_757
timestamp 1636968456
transform 1 0 71668 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_769
timestamp 1636968456
transform 1 0 72772 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_781
timestamp 1636968456
transform 1 0 73876 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_793
timestamp 1636968456
transform 1 0 74980 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_805
timestamp 1
transform 1 0 76084 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_811
timestamp 1
transform 1 0 76636 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_813
timestamp 1
transform 1 0 76820 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_128_821
timestamp 1
transform 1 0 77556 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_3
timestamp 1636968456
transform 1 0 2300 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_15
timestamp 1636968456
transform 1 0 3404 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_27
timestamp 1636968456
transform 1 0 4508 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_39
timestamp 1636968456
transform 1 0 5612 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_129_51
timestamp 1
transform 1 0 6716 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1
transform 1 0 7084 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_57
timestamp 1636968456
transform 1 0 7268 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_69
timestamp 1636968456
transform 1 0 8372 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_81
timestamp 1636968456
transform 1 0 9476 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_93
timestamp 1636968456
transform 1 0 10580 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_105
timestamp 1
transform 1 0 11684 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_111
timestamp 1
transform 1 0 12236 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_113
timestamp 1636968456
transform 1 0 12420 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_125
timestamp 1636968456
transform 1 0 13524 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_137
timestamp 1636968456
transform 1 0 14628 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_149
timestamp 1636968456
transform 1 0 15732 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_161
timestamp 1
transform 1 0 16836 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_167
timestamp 1
transform 1 0 17388 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_169
timestamp 1636968456
transform 1 0 17572 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_181
timestamp 1636968456
transform 1 0 18676 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_193
timestamp 1636968456
transform 1 0 19780 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_205
timestamp 1636968456
transform 1 0 20884 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_217
timestamp 1
transform 1 0 21988 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_223
timestamp 1
transform 1 0 22540 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_225
timestamp 1636968456
transform 1 0 22724 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_237
timestamp 1636968456
transform 1 0 23828 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_249
timestamp 1636968456
transform 1 0 24932 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_261
timestamp 1636968456
transform 1 0 26036 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_273
timestamp 1
transform 1 0 27140 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_279
timestamp 1
transform 1 0 27692 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_281
timestamp 1636968456
transform 1 0 27876 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_293
timestamp 1636968456
transform 1 0 28980 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_305
timestamp 1636968456
transform 1 0 30084 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_317
timestamp 1636968456
transform 1 0 31188 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_329
timestamp 1
transform 1 0 32292 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_335
timestamp 1
transform 1 0 32844 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_337
timestamp 1636968456
transform 1 0 33028 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_349
timestamp 1636968456
transform 1 0 34132 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_361
timestamp 1636968456
transform 1 0 35236 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_373
timestamp 1636968456
transform 1 0 36340 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_385
timestamp 1
transform 1 0 37444 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_391
timestamp 1
transform 1 0 37996 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_393
timestamp 1636968456
transform 1 0 38180 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_405
timestamp 1636968456
transform 1 0 39284 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_417
timestamp 1636968456
transform 1 0 40388 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_429
timestamp 1636968456
transform 1 0 41492 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_441
timestamp 1
transform 1 0 42596 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_447
timestamp 1
transform 1 0 43148 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_449
timestamp 1636968456
transform 1 0 43332 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_461
timestamp 1636968456
transform 1 0 44436 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_473
timestamp 1636968456
transform 1 0 45540 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_485
timestamp 1636968456
transform 1 0 46644 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_497
timestamp 1
transform 1 0 47748 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_503
timestamp 1
transform 1 0 48300 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_505
timestamp 1636968456
transform 1 0 48484 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_517
timestamp 1636968456
transform 1 0 49588 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_529
timestamp 1636968456
transform 1 0 50692 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_541
timestamp 1636968456
transform 1 0 51796 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_553
timestamp 1
transform 1 0 52900 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_559
timestamp 1
transform 1 0 53452 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_561
timestamp 1636968456
transform 1 0 53636 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_573
timestamp 1636968456
transform 1 0 54740 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_585
timestamp 1636968456
transform 1 0 55844 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_597
timestamp 1636968456
transform 1 0 56948 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_609
timestamp 1
transform 1 0 58052 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_615
timestamp 1
transform 1 0 58604 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_617
timestamp 1636968456
transform 1 0 58788 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_629
timestamp 1636968456
transform 1 0 59892 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_641
timestamp 1636968456
transform 1 0 60996 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_653
timestamp 1636968456
transform 1 0 62100 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_665
timestamp 1
transform 1 0 63204 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_671
timestamp 1
transform 1 0 63756 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_673
timestamp 1636968456
transform 1 0 63940 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_685
timestamp 1636968456
transform 1 0 65044 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_697
timestamp 1636968456
transform 1 0 66148 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_709
timestamp 1636968456
transform 1 0 67252 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_721
timestamp 1
transform 1 0 68356 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_727
timestamp 1
transform 1 0 68908 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_729
timestamp 1636968456
transform 1 0 69092 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_741
timestamp 1636968456
transform 1 0 70196 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_753
timestamp 1636968456
transform 1 0 71300 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_765
timestamp 1636968456
transform 1 0 72404 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_777
timestamp 1
transform 1 0 73508 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_783
timestamp 1
transform 1 0 74060 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_785
timestamp 1636968456
transform 1 0 74244 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_797
timestamp 1636968456
transform 1 0 75348 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_809
timestamp 1636968456
transform 1 0 76452 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_129_821
timestamp 1
transform 1 0 77556 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_3
timestamp 1636968456
transform 1 0 2300 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_15
timestamp 1636968456
transform 1 0 3404 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 1
transform 1 0 4508 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_29
timestamp 1636968456
transform 1 0 4692 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_41
timestamp 1636968456
transform 1 0 5796 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_53
timestamp 1636968456
transform 1 0 6900 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_65
timestamp 1636968456
transform 1 0 8004 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1
transform 1 0 9108 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1
transform 1 0 9660 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_85
timestamp 1636968456
transform 1 0 9844 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_97
timestamp 1636968456
transform 1 0 10948 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_109
timestamp 1636968456
transform 1 0 12052 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_121
timestamp 1636968456
transform 1 0 13156 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_133
timestamp 1
transform 1 0 14260 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_139
timestamp 1
transform 1 0 14812 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_141
timestamp 1636968456
transform 1 0 14996 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_153
timestamp 1636968456
transform 1 0 16100 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_165
timestamp 1636968456
transform 1 0 17204 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_177
timestamp 1636968456
transform 1 0 18308 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_189
timestamp 1
transform 1 0 19412 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_195
timestamp 1
transform 1 0 19964 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_197
timestamp 1636968456
transform 1 0 20148 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_209
timestamp 1636968456
transform 1 0 21252 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_221
timestamp 1636968456
transform 1 0 22356 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_233
timestamp 1636968456
transform 1 0 23460 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_245
timestamp 1
transform 1 0 24564 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_251
timestamp 1
transform 1 0 25116 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_253
timestamp 1636968456
transform 1 0 25300 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_265
timestamp 1636968456
transform 1 0 26404 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_277
timestamp 1636968456
transform 1 0 27508 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_289
timestamp 1636968456
transform 1 0 28612 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_301
timestamp 1
transform 1 0 29716 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_307
timestamp 1
transform 1 0 30268 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_309
timestamp 1636968456
transform 1 0 30452 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_321
timestamp 1636968456
transform 1 0 31556 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_333
timestamp 1636968456
transform 1 0 32660 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_345
timestamp 1636968456
transform 1 0 33764 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_357
timestamp 1
transform 1 0 34868 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_363
timestamp 1
transform 1 0 35420 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_365
timestamp 1636968456
transform 1 0 35604 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_377
timestamp 1636968456
transform 1 0 36708 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_389
timestamp 1636968456
transform 1 0 37812 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_401
timestamp 1636968456
transform 1 0 38916 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_413
timestamp 1
transform 1 0 40020 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_419
timestamp 1
transform 1 0 40572 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_421
timestamp 1636968456
transform 1 0 40756 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_433
timestamp 1636968456
transform 1 0 41860 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_445
timestamp 1636968456
transform 1 0 42964 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_457
timestamp 1636968456
transform 1 0 44068 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_469
timestamp 1
transform 1 0 45172 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_475
timestamp 1
transform 1 0 45724 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_477
timestamp 1636968456
transform 1 0 45908 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_489
timestamp 1636968456
transform 1 0 47012 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_501
timestamp 1636968456
transform 1 0 48116 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_513
timestamp 1636968456
transform 1 0 49220 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_525
timestamp 1
transform 1 0 50324 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_531
timestamp 1
transform 1 0 50876 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_533
timestamp 1636968456
transform 1 0 51060 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_545
timestamp 1636968456
transform 1 0 52164 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_557
timestamp 1636968456
transform 1 0 53268 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_569
timestamp 1636968456
transform 1 0 54372 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_581
timestamp 1
transform 1 0 55476 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_587
timestamp 1
transform 1 0 56028 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_589
timestamp 1636968456
transform 1 0 56212 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_601
timestamp 1636968456
transform 1 0 57316 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_613
timestamp 1636968456
transform 1 0 58420 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_625
timestamp 1636968456
transform 1 0 59524 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_637
timestamp 1
transform 1 0 60628 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_643
timestamp 1
transform 1 0 61180 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_645
timestamp 1636968456
transform 1 0 61364 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_657
timestamp 1636968456
transform 1 0 62468 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_669
timestamp 1636968456
transform 1 0 63572 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_681
timestamp 1636968456
transform 1 0 64676 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_693
timestamp 1
transform 1 0 65780 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_699
timestamp 1
transform 1 0 66332 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_701
timestamp 1636968456
transform 1 0 66516 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_713
timestamp 1636968456
transform 1 0 67620 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_725
timestamp 1636968456
transform 1 0 68724 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_737
timestamp 1636968456
transform 1 0 69828 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_749
timestamp 1
transform 1 0 70932 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_755
timestamp 1
transform 1 0 71484 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_757
timestamp 1636968456
transform 1 0 71668 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_769
timestamp 1636968456
transform 1 0 72772 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_781
timestamp 1636968456
transform 1 0 73876 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_793
timestamp 1636968456
transform 1 0 74980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_805
timestamp 1
transform 1 0 76084 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_811
timestamp 1
transform 1 0 76636 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_813
timestamp 1
transform 1 0 76820 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_821
timestamp 1
transform 1 0 77556 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_3
timestamp 1636968456
transform 1 0 2300 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_15
timestamp 1636968456
transform 1 0 3404 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_27
timestamp 1636968456
transform 1 0 4508 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_39
timestamp 1636968456
transform 1 0 5612 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_51
timestamp 1
transform 1 0 6716 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_55
timestamp 1
transform 1 0 7084 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_57
timestamp 1636968456
transform 1 0 7268 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_69
timestamp 1636968456
transform 1 0 8372 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_81
timestamp 1636968456
transform 1 0 9476 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_93
timestamp 1636968456
transform 1 0 10580 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_105
timestamp 1
transform 1 0 11684 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_111
timestamp 1
transform 1 0 12236 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_113
timestamp 1636968456
transform 1 0 12420 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_125
timestamp 1636968456
transform 1 0 13524 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_137
timestamp 1636968456
transform 1 0 14628 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_149
timestamp 1636968456
transform 1 0 15732 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_161
timestamp 1
transform 1 0 16836 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_167
timestamp 1
transform 1 0 17388 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_169
timestamp 1636968456
transform 1 0 17572 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_181
timestamp 1636968456
transform 1 0 18676 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_193
timestamp 1636968456
transform 1 0 19780 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_205
timestamp 1636968456
transform 1 0 20884 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_217
timestamp 1
transform 1 0 21988 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_223
timestamp 1
transform 1 0 22540 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_225
timestamp 1636968456
transform 1 0 22724 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_237
timestamp 1636968456
transform 1 0 23828 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_249
timestamp 1636968456
transform 1 0 24932 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_261
timestamp 1636968456
transform 1 0 26036 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_273
timestamp 1
transform 1 0 27140 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_279
timestamp 1
transform 1 0 27692 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_281
timestamp 1636968456
transform 1 0 27876 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_293
timestamp 1636968456
transform 1 0 28980 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_305
timestamp 1636968456
transform 1 0 30084 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_317
timestamp 1636968456
transform 1 0 31188 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_329
timestamp 1
transform 1 0 32292 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_335
timestamp 1
transform 1 0 32844 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_337
timestamp 1636968456
transform 1 0 33028 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_349
timestamp 1636968456
transform 1 0 34132 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_361
timestamp 1636968456
transform 1 0 35236 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_373
timestamp 1636968456
transform 1 0 36340 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_385
timestamp 1
transform 1 0 37444 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_391
timestamp 1
transform 1 0 37996 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_393
timestamp 1636968456
transform 1 0 38180 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_405
timestamp 1636968456
transform 1 0 39284 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_417
timestamp 1636968456
transform 1 0 40388 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_429
timestamp 1636968456
transform 1 0 41492 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_441
timestamp 1
transform 1 0 42596 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_447
timestamp 1
transform 1 0 43148 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_449
timestamp 1636968456
transform 1 0 43332 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_461
timestamp 1636968456
transform 1 0 44436 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_473
timestamp 1636968456
transform 1 0 45540 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_485
timestamp 1636968456
transform 1 0 46644 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_497
timestamp 1
transform 1 0 47748 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_503
timestamp 1
transform 1 0 48300 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_505
timestamp 1636968456
transform 1 0 48484 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_517
timestamp 1636968456
transform 1 0 49588 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_529
timestamp 1636968456
transform 1 0 50692 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_541
timestamp 1636968456
transform 1 0 51796 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_553
timestamp 1
transform 1 0 52900 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_559
timestamp 1
transform 1 0 53452 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_561
timestamp 1636968456
transform 1 0 53636 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_573
timestamp 1636968456
transform 1 0 54740 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_585
timestamp 1636968456
transform 1 0 55844 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_597
timestamp 1636968456
transform 1 0 56948 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_609
timestamp 1
transform 1 0 58052 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_615
timestamp 1
transform 1 0 58604 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_617
timestamp 1636968456
transform 1 0 58788 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_629
timestamp 1636968456
transform 1 0 59892 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_641
timestamp 1636968456
transform 1 0 60996 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_653
timestamp 1636968456
transform 1 0 62100 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_665
timestamp 1
transform 1 0 63204 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_671
timestamp 1
transform 1 0 63756 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_673
timestamp 1636968456
transform 1 0 63940 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_685
timestamp 1636968456
transform 1 0 65044 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_697
timestamp 1636968456
transform 1 0 66148 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_709
timestamp 1636968456
transform 1 0 67252 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_721
timestamp 1
transform 1 0 68356 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_727
timestamp 1
transform 1 0 68908 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_729
timestamp 1636968456
transform 1 0 69092 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_741
timestamp 1636968456
transform 1 0 70196 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_753
timestamp 1636968456
transform 1 0 71300 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_765
timestamp 1636968456
transform 1 0 72404 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_777
timestamp 1
transform 1 0 73508 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_783
timestamp 1
transform 1 0 74060 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_785
timestamp 1636968456
transform 1 0 74244 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_797
timestamp 1636968456
transform 1 0 75348 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_809
timestamp 1636968456
transform 1 0 76452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_131_821
timestamp 1
transform 1 0 77556 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_3
timestamp 1636968456
transform 1 0 2300 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_15
timestamp 1636968456
transform 1 0 3404 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1
transform 1 0 4508 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_29
timestamp 1636968456
transform 1 0 4692 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_41
timestamp 1636968456
transform 1 0 5796 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_53
timestamp 1636968456
transform 1 0 6900 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_65
timestamp 1636968456
transform 1 0 8004 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1
transform 1 0 9108 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1
transform 1 0 9660 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_85
timestamp 1636968456
transform 1 0 9844 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_97
timestamp 1636968456
transform 1 0 10948 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_109
timestamp 1636968456
transform 1 0 12052 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_121
timestamp 1636968456
transform 1 0 13156 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_133
timestamp 1
transform 1 0 14260 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_139
timestamp 1
transform 1 0 14812 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_141
timestamp 1636968456
transform 1 0 14996 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_153
timestamp 1636968456
transform 1 0 16100 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_165
timestamp 1636968456
transform 1 0 17204 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_177
timestamp 1636968456
transform 1 0 18308 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_189
timestamp 1
transform 1 0 19412 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_195
timestamp 1
transform 1 0 19964 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_197
timestamp 1636968456
transform 1 0 20148 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_209
timestamp 1636968456
transform 1 0 21252 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_221
timestamp 1636968456
transform 1 0 22356 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_233
timestamp 1636968456
transform 1 0 23460 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_245
timestamp 1
transform 1 0 24564 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_251
timestamp 1
transform 1 0 25116 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_253
timestamp 1636968456
transform 1 0 25300 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_265
timestamp 1636968456
transform 1 0 26404 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_277
timestamp 1636968456
transform 1 0 27508 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_289
timestamp 1636968456
transform 1 0 28612 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_301
timestamp 1
transform 1 0 29716 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_307
timestamp 1
transform 1 0 30268 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_309
timestamp 1636968456
transform 1 0 30452 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_321
timestamp 1636968456
transform 1 0 31556 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_333
timestamp 1636968456
transform 1 0 32660 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_345
timestamp 1636968456
transform 1 0 33764 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_357
timestamp 1
transform 1 0 34868 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_363
timestamp 1
transform 1 0 35420 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_365
timestamp 1636968456
transform 1 0 35604 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_377
timestamp 1636968456
transform 1 0 36708 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_389
timestamp 1636968456
transform 1 0 37812 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_401
timestamp 1636968456
transform 1 0 38916 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_413
timestamp 1
transform 1 0 40020 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_419
timestamp 1
transform 1 0 40572 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_421
timestamp 1636968456
transform 1 0 40756 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_433
timestamp 1636968456
transform 1 0 41860 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_445
timestamp 1636968456
transform 1 0 42964 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_457
timestamp 1636968456
transform 1 0 44068 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_469
timestamp 1
transform 1 0 45172 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_475
timestamp 1
transform 1 0 45724 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_477
timestamp 1636968456
transform 1 0 45908 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_489
timestamp 1636968456
transform 1 0 47012 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_501
timestamp 1636968456
transform 1 0 48116 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_513
timestamp 1636968456
transform 1 0 49220 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_525
timestamp 1
transform 1 0 50324 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_531
timestamp 1
transform 1 0 50876 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_533
timestamp 1636968456
transform 1 0 51060 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_545
timestamp 1636968456
transform 1 0 52164 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_557
timestamp 1636968456
transform 1 0 53268 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_569
timestamp 1636968456
transform 1 0 54372 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_581
timestamp 1
transform 1 0 55476 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_587
timestamp 1
transform 1 0 56028 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_589
timestamp 1636968456
transform 1 0 56212 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_601
timestamp 1636968456
transform 1 0 57316 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_613
timestamp 1636968456
transform 1 0 58420 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_625
timestamp 1636968456
transform 1 0 59524 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_637
timestamp 1
transform 1 0 60628 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_643
timestamp 1
transform 1 0 61180 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_645
timestamp 1636968456
transform 1 0 61364 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_657
timestamp 1636968456
transform 1 0 62468 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_669
timestamp 1636968456
transform 1 0 63572 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_681
timestamp 1636968456
transform 1 0 64676 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_693
timestamp 1
transform 1 0 65780 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_699
timestamp 1
transform 1 0 66332 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_701
timestamp 1636968456
transform 1 0 66516 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_713
timestamp 1636968456
transform 1 0 67620 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_725
timestamp 1636968456
transform 1 0 68724 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_737
timestamp 1636968456
transform 1 0 69828 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_749
timestamp 1
transform 1 0 70932 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_755
timestamp 1
transform 1 0 71484 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_757
timestamp 1636968456
transform 1 0 71668 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_769
timestamp 1636968456
transform 1 0 72772 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_781
timestamp 1636968456
transform 1 0 73876 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_793
timestamp 1636968456
transform 1 0 74980 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_805
timestamp 1
transform 1 0 76084 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_811
timestamp 1
transform 1 0 76636 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_813
timestamp 1
transform 1 0 76820 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_821
timestamp 1
transform 1 0 77556 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1636968456
transform 1 0 2300 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1636968456
transform 1 0 3404 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_27
timestamp 1636968456
transform 1 0 4508 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_39
timestamp 1636968456
transform 1 0 5612 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_51
timestamp 1
transform 1 0 6716 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_55
timestamp 1
transform 1 0 7084 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_57
timestamp 1636968456
transform 1 0 7268 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_69
timestamp 1636968456
transform 1 0 8372 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_81
timestamp 1636968456
transform 1 0 9476 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_93
timestamp 1636968456
transform 1 0 10580 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_105
timestamp 1
transform 1 0 11684 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_111
timestamp 1
transform 1 0 12236 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_113
timestamp 1636968456
transform 1 0 12420 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_125
timestamp 1636968456
transform 1 0 13524 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_137
timestamp 1636968456
transform 1 0 14628 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_149
timestamp 1636968456
transform 1 0 15732 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_161
timestamp 1
transform 1 0 16836 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_167
timestamp 1
transform 1 0 17388 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_169
timestamp 1636968456
transform 1 0 17572 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_181
timestamp 1636968456
transform 1 0 18676 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_193
timestamp 1636968456
transform 1 0 19780 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_205
timestamp 1636968456
transform 1 0 20884 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_217
timestamp 1
transform 1 0 21988 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_223
timestamp 1
transform 1 0 22540 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_225
timestamp 1636968456
transform 1 0 22724 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_237
timestamp 1636968456
transform 1 0 23828 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_249
timestamp 1636968456
transform 1 0 24932 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_261
timestamp 1636968456
transform 1 0 26036 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_273
timestamp 1
transform 1 0 27140 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_279
timestamp 1
transform 1 0 27692 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_281
timestamp 1636968456
transform 1 0 27876 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_293
timestamp 1636968456
transform 1 0 28980 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_305
timestamp 1636968456
transform 1 0 30084 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_317
timestamp 1636968456
transform 1 0 31188 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_329
timestamp 1
transform 1 0 32292 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_335
timestamp 1
transform 1 0 32844 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_337
timestamp 1636968456
transform 1 0 33028 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_349
timestamp 1636968456
transform 1 0 34132 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_361
timestamp 1636968456
transform 1 0 35236 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_373
timestamp 1636968456
transform 1 0 36340 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_385
timestamp 1
transform 1 0 37444 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_391
timestamp 1
transform 1 0 37996 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_393
timestamp 1636968456
transform 1 0 38180 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_405
timestamp 1636968456
transform 1 0 39284 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_417
timestamp 1636968456
transform 1 0 40388 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_429
timestamp 1636968456
transform 1 0 41492 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_441
timestamp 1
transform 1 0 42596 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_447
timestamp 1
transform 1 0 43148 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_449
timestamp 1636968456
transform 1 0 43332 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_461
timestamp 1636968456
transform 1 0 44436 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_473
timestamp 1636968456
transform 1 0 45540 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_485
timestamp 1636968456
transform 1 0 46644 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_497
timestamp 1
transform 1 0 47748 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_503
timestamp 1
transform 1 0 48300 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_505
timestamp 1636968456
transform 1 0 48484 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_517
timestamp 1636968456
transform 1 0 49588 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_529
timestamp 1636968456
transform 1 0 50692 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_541
timestamp 1636968456
transform 1 0 51796 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_553
timestamp 1
transform 1 0 52900 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_559
timestamp 1
transform 1 0 53452 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_561
timestamp 1636968456
transform 1 0 53636 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_573
timestamp 1636968456
transform 1 0 54740 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_585
timestamp 1636968456
transform 1 0 55844 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_597
timestamp 1636968456
transform 1 0 56948 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_609
timestamp 1
transform 1 0 58052 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_615
timestamp 1
transform 1 0 58604 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_617
timestamp 1636968456
transform 1 0 58788 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_629
timestamp 1636968456
transform 1 0 59892 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_641
timestamp 1636968456
transform 1 0 60996 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_653
timestamp 1636968456
transform 1 0 62100 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_665
timestamp 1
transform 1 0 63204 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_671
timestamp 1
transform 1 0 63756 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_673
timestamp 1636968456
transform 1 0 63940 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_685
timestamp 1636968456
transform 1 0 65044 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_697
timestamp 1636968456
transform 1 0 66148 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_709
timestamp 1636968456
transform 1 0 67252 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_721
timestamp 1
transform 1 0 68356 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_727
timestamp 1
transform 1 0 68908 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_729
timestamp 1636968456
transform 1 0 69092 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_741
timestamp 1636968456
transform 1 0 70196 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_753
timestamp 1636968456
transform 1 0 71300 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_765
timestamp 1636968456
transform 1 0 72404 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_777
timestamp 1
transform 1 0 73508 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_783
timestamp 1
transform 1 0 74060 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_785
timestamp 1636968456
transform 1 0 74244 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_797
timestamp 1636968456
transform 1 0 75348 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_809
timestamp 1636968456
transform 1 0 76452 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_133_821
timestamp 1
transform 1 0 77556 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_3
timestamp 1636968456
transform 1 0 2300 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_15
timestamp 1636968456
transform 1 0 3404 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1
transform 1 0 4508 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_29
timestamp 1636968456
transform 1 0 4692 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_41
timestamp 1636968456
transform 1 0 5796 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_53
timestamp 1636968456
transform 1 0 6900 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_65
timestamp 1636968456
transform 1 0 8004 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1
transform 1 0 9108 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1
transform 1 0 9660 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_85
timestamp 1636968456
transform 1 0 9844 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_97
timestamp 1636968456
transform 1 0 10948 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_109
timestamp 1636968456
transform 1 0 12052 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_121
timestamp 1636968456
transform 1 0 13156 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_133
timestamp 1
transform 1 0 14260 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_139
timestamp 1
transform 1 0 14812 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_141
timestamp 1636968456
transform 1 0 14996 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_153
timestamp 1636968456
transform 1 0 16100 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_165
timestamp 1636968456
transform 1 0 17204 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_177
timestamp 1636968456
transform 1 0 18308 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_189
timestamp 1
transform 1 0 19412 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_195
timestamp 1
transform 1 0 19964 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_197
timestamp 1636968456
transform 1 0 20148 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_209
timestamp 1636968456
transform 1 0 21252 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_221
timestamp 1636968456
transform 1 0 22356 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_233
timestamp 1636968456
transform 1 0 23460 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_245
timestamp 1
transform 1 0 24564 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_251
timestamp 1
transform 1 0 25116 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_253
timestamp 1636968456
transform 1 0 25300 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_265
timestamp 1636968456
transform 1 0 26404 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_277
timestamp 1636968456
transform 1 0 27508 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_289
timestamp 1636968456
transform 1 0 28612 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_301
timestamp 1
transform 1 0 29716 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_307
timestamp 1
transform 1 0 30268 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_309
timestamp 1636968456
transform 1 0 30452 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_321
timestamp 1636968456
transform 1 0 31556 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_333
timestamp 1636968456
transform 1 0 32660 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_345
timestamp 1636968456
transform 1 0 33764 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_357
timestamp 1
transform 1 0 34868 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_363
timestamp 1
transform 1 0 35420 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_365
timestamp 1636968456
transform 1 0 35604 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_377
timestamp 1636968456
transform 1 0 36708 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_389
timestamp 1636968456
transform 1 0 37812 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_401
timestamp 1636968456
transform 1 0 38916 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_413
timestamp 1
transform 1 0 40020 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_419
timestamp 1
transform 1 0 40572 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_421
timestamp 1636968456
transform 1 0 40756 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_433
timestamp 1636968456
transform 1 0 41860 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_445
timestamp 1636968456
transform 1 0 42964 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_457
timestamp 1636968456
transform 1 0 44068 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_469
timestamp 1
transform 1 0 45172 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_475
timestamp 1
transform 1 0 45724 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_477
timestamp 1636968456
transform 1 0 45908 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_489
timestamp 1636968456
transform 1 0 47012 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_501
timestamp 1636968456
transform 1 0 48116 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_513
timestamp 1636968456
transform 1 0 49220 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_525
timestamp 1
transform 1 0 50324 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_531
timestamp 1
transform 1 0 50876 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_533
timestamp 1636968456
transform 1 0 51060 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_545
timestamp 1636968456
transform 1 0 52164 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_557
timestamp 1636968456
transform 1 0 53268 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_569
timestamp 1636968456
transform 1 0 54372 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_581
timestamp 1
transform 1 0 55476 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_587
timestamp 1
transform 1 0 56028 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_589
timestamp 1636968456
transform 1 0 56212 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_601
timestamp 1636968456
transform 1 0 57316 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_613
timestamp 1636968456
transform 1 0 58420 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_625
timestamp 1636968456
transform 1 0 59524 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_637
timestamp 1
transform 1 0 60628 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_643
timestamp 1
transform 1 0 61180 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_645
timestamp 1636968456
transform 1 0 61364 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_657
timestamp 1636968456
transform 1 0 62468 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_669
timestamp 1636968456
transform 1 0 63572 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_681
timestamp 1636968456
transform 1 0 64676 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_693
timestamp 1
transform 1 0 65780 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_699
timestamp 1
transform 1 0 66332 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_701
timestamp 1636968456
transform 1 0 66516 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_713
timestamp 1636968456
transform 1 0 67620 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_725
timestamp 1636968456
transform 1 0 68724 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_737
timestamp 1636968456
transform 1 0 69828 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_749
timestamp 1
transform 1 0 70932 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_755
timestamp 1
transform 1 0 71484 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_757
timestamp 1636968456
transform 1 0 71668 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_769
timestamp 1636968456
transform 1 0 72772 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_781
timestamp 1636968456
transform 1 0 73876 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_793
timestamp 1636968456
transform 1 0 74980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_805
timestamp 1
transform 1 0 76084 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_811
timestamp 1
transform 1 0 76636 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_813
timestamp 1
transform 1 0 76820 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_821
timestamp 1
transform 1 0 77556 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_3
timestamp 1636968456
transform 1 0 2300 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_15
timestamp 1636968456
transform 1 0 3404 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_27
timestamp 1636968456
transform 1 0 4508 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_39
timestamp 1636968456
transform 1 0 5612 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_51
timestamp 1
transform 1 0 6716 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_55
timestamp 1
transform 1 0 7084 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_57
timestamp 1636968456
transform 1 0 7268 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_69
timestamp 1636968456
transform 1 0 8372 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_81
timestamp 1636968456
transform 1 0 9476 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_93
timestamp 1636968456
transform 1 0 10580 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_105
timestamp 1
transform 1 0 11684 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_111
timestamp 1
transform 1 0 12236 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_113
timestamp 1636968456
transform 1 0 12420 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_125
timestamp 1636968456
transform 1 0 13524 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_137
timestamp 1636968456
transform 1 0 14628 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_149
timestamp 1636968456
transform 1 0 15732 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_161
timestamp 1
transform 1 0 16836 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_167
timestamp 1
transform 1 0 17388 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_169
timestamp 1636968456
transform 1 0 17572 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_181
timestamp 1636968456
transform 1 0 18676 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_193
timestamp 1636968456
transform 1 0 19780 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_205
timestamp 1636968456
transform 1 0 20884 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_217
timestamp 1
transform 1 0 21988 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_223
timestamp 1
transform 1 0 22540 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_225
timestamp 1636968456
transform 1 0 22724 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_237
timestamp 1636968456
transform 1 0 23828 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_249
timestamp 1636968456
transform 1 0 24932 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_261
timestamp 1636968456
transform 1 0 26036 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_273
timestamp 1
transform 1 0 27140 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_279
timestamp 1
transform 1 0 27692 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_281
timestamp 1636968456
transform 1 0 27876 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_293
timestamp 1636968456
transform 1 0 28980 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_305
timestamp 1636968456
transform 1 0 30084 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_317
timestamp 1636968456
transform 1 0 31188 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_329
timestamp 1
transform 1 0 32292 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_335
timestamp 1
transform 1 0 32844 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_337
timestamp 1636968456
transform 1 0 33028 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_349
timestamp 1636968456
transform 1 0 34132 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_361
timestamp 1636968456
transform 1 0 35236 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_373
timestamp 1636968456
transform 1 0 36340 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_385
timestamp 1
transform 1 0 37444 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_391
timestamp 1
transform 1 0 37996 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_393
timestamp 1636968456
transform 1 0 38180 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_405
timestamp 1636968456
transform 1 0 39284 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_417
timestamp 1636968456
transform 1 0 40388 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_429
timestamp 1636968456
transform 1 0 41492 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_441
timestamp 1
transform 1 0 42596 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_447
timestamp 1
transform 1 0 43148 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_449
timestamp 1636968456
transform 1 0 43332 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_461
timestamp 1636968456
transform 1 0 44436 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_473
timestamp 1636968456
transform 1 0 45540 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_485
timestamp 1636968456
transform 1 0 46644 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_497
timestamp 1
transform 1 0 47748 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_503
timestamp 1
transform 1 0 48300 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_505
timestamp 1636968456
transform 1 0 48484 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_517
timestamp 1636968456
transform 1 0 49588 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_529
timestamp 1636968456
transform 1 0 50692 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_541
timestamp 1636968456
transform 1 0 51796 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_553
timestamp 1
transform 1 0 52900 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_559
timestamp 1
transform 1 0 53452 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_561
timestamp 1636968456
transform 1 0 53636 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_573
timestamp 1636968456
transform 1 0 54740 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_585
timestamp 1636968456
transform 1 0 55844 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_597
timestamp 1636968456
transform 1 0 56948 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_609
timestamp 1
transform 1 0 58052 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_615
timestamp 1
transform 1 0 58604 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_617
timestamp 1636968456
transform 1 0 58788 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_629
timestamp 1636968456
transform 1 0 59892 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_641
timestamp 1636968456
transform 1 0 60996 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_653
timestamp 1636968456
transform 1 0 62100 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_665
timestamp 1
transform 1 0 63204 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_671
timestamp 1
transform 1 0 63756 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_673
timestamp 1636968456
transform 1 0 63940 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_685
timestamp 1636968456
transform 1 0 65044 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_697
timestamp 1636968456
transform 1 0 66148 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_709
timestamp 1636968456
transform 1 0 67252 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_721
timestamp 1
transform 1 0 68356 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_727
timestamp 1
transform 1 0 68908 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_729
timestamp 1636968456
transform 1 0 69092 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_741
timestamp 1636968456
transform 1 0 70196 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_753
timestamp 1636968456
transform 1 0 71300 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_765
timestamp 1636968456
transform 1 0 72404 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_777
timestamp 1
transform 1 0 73508 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_783
timestamp 1
transform 1 0 74060 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_785
timestamp 1636968456
transform 1 0 74244 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_797
timestamp 1636968456
transform 1 0 75348 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_809
timestamp 1636968456
transform 1 0 76452 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_135_821
timestamp 1
transform 1 0 77556 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_3
timestamp 1636968456
transform 1 0 2300 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_15
timestamp 1636968456
transform 1 0 3404 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1
transform 1 0 4508 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_29
timestamp 1636968456
transform 1 0 4692 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_41
timestamp 1636968456
transform 1 0 5796 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_53
timestamp 1636968456
transform 1 0 6900 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_65
timestamp 1636968456
transform 1 0 8004 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1
transform 1 0 9108 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1
transform 1 0 9660 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_85
timestamp 1636968456
transform 1 0 9844 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_97
timestamp 1636968456
transform 1 0 10948 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_109
timestamp 1636968456
transform 1 0 12052 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_121
timestamp 1636968456
transform 1 0 13156 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_133
timestamp 1
transform 1 0 14260 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_139
timestamp 1
transform 1 0 14812 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_141
timestamp 1636968456
transform 1 0 14996 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_153
timestamp 1636968456
transform 1 0 16100 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_165
timestamp 1636968456
transform 1 0 17204 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_177
timestamp 1636968456
transform 1 0 18308 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_189
timestamp 1
transform 1 0 19412 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_195
timestamp 1
transform 1 0 19964 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_197
timestamp 1636968456
transform 1 0 20148 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_209
timestamp 1636968456
transform 1 0 21252 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_221
timestamp 1636968456
transform 1 0 22356 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_233
timestamp 1636968456
transform 1 0 23460 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_245
timestamp 1
transform 1 0 24564 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_251
timestamp 1
transform 1 0 25116 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_253
timestamp 1636968456
transform 1 0 25300 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_265
timestamp 1636968456
transform 1 0 26404 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_277
timestamp 1636968456
transform 1 0 27508 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_289
timestamp 1636968456
transform 1 0 28612 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_301
timestamp 1
transform 1 0 29716 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_307
timestamp 1
transform 1 0 30268 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_309
timestamp 1636968456
transform 1 0 30452 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_321
timestamp 1636968456
transform 1 0 31556 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_333
timestamp 1636968456
transform 1 0 32660 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_345
timestamp 1636968456
transform 1 0 33764 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_357
timestamp 1
transform 1 0 34868 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_363
timestamp 1
transform 1 0 35420 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_365
timestamp 1636968456
transform 1 0 35604 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_377
timestamp 1636968456
transform 1 0 36708 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_389
timestamp 1636968456
transform 1 0 37812 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_401
timestamp 1636968456
transform 1 0 38916 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_413
timestamp 1
transform 1 0 40020 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_419
timestamp 1
transform 1 0 40572 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_421
timestamp 1636968456
transform 1 0 40756 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_433
timestamp 1636968456
transform 1 0 41860 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_445
timestamp 1636968456
transform 1 0 42964 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_457
timestamp 1636968456
transform 1 0 44068 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_469
timestamp 1
transform 1 0 45172 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_475
timestamp 1
transform 1 0 45724 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_477
timestamp 1636968456
transform 1 0 45908 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_489
timestamp 1636968456
transform 1 0 47012 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_501
timestamp 1636968456
transform 1 0 48116 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_513
timestamp 1636968456
transform 1 0 49220 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_525
timestamp 1
transform 1 0 50324 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_531
timestamp 1
transform 1 0 50876 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_533
timestamp 1636968456
transform 1 0 51060 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_545
timestamp 1636968456
transform 1 0 52164 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_557
timestamp 1636968456
transform 1 0 53268 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_569
timestamp 1636968456
transform 1 0 54372 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_581
timestamp 1
transform 1 0 55476 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_587
timestamp 1
transform 1 0 56028 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_589
timestamp 1636968456
transform 1 0 56212 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_601
timestamp 1636968456
transform 1 0 57316 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_613
timestamp 1636968456
transform 1 0 58420 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_625
timestamp 1636968456
transform 1 0 59524 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_637
timestamp 1
transform 1 0 60628 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_643
timestamp 1
transform 1 0 61180 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_645
timestamp 1636968456
transform 1 0 61364 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_657
timestamp 1636968456
transform 1 0 62468 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_669
timestamp 1636968456
transform 1 0 63572 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_681
timestamp 1636968456
transform 1 0 64676 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_693
timestamp 1
transform 1 0 65780 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_699
timestamp 1
transform 1 0 66332 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_701
timestamp 1636968456
transform 1 0 66516 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_713
timestamp 1636968456
transform 1 0 67620 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_725
timestamp 1636968456
transform 1 0 68724 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_737
timestamp 1636968456
transform 1 0 69828 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_749
timestamp 1
transform 1 0 70932 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_755
timestamp 1
transform 1 0 71484 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_757
timestamp 1636968456
transform 1 0 71668 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_769
timestamp 1636968456
transform 1 0 72772 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_781
timestamp 1636968456
transform 1 0 73876 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_793
timestamp 1636968456
transform 1 0 74980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_805
timestamp 1
transform 1 0 76084 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_811
timestamp 1
transform 1 0 76636 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_813
timestamp 1
transform 1 0 76820 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_821
timestamp 1
transform 1 0 77556 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_3
timestamp 1636968456
transform 1 0 2300 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_15
timestamp 1636968456
transform 1 0 3404 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_27
timestamp 1636968456
transform 1 0 4508 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_39
timestamp 1636968456
transform 1 0 5612 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_51
timestamp 1
transform 1 0 6716 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1
transform 1 0 7084 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_57
timestamp 1636968456
transform 1 0 7268 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_69
timestamp 1636968456
transform 1 0 8372 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_81
timestamp 1636968456
transform 1 0 9476 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_93
timestamp 1636968456
transform 1 0 10580 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_105
timestamp 1
transform 1 0 11684 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_111
timestamp 1
transform 1 0 12236 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_113
timestamp 1636968456
transform 1 0 12420 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_125
timestamp 1636968456
transform 1 0 13524 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_137
timestamp 1636968456
transform 1 0 14628 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_149
timestamp 1636968456
transform 1 0 15732 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_161
timestamp 1
transform 1 0 16836 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_167
timestamp 1
transform 1 0 17388 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_169
timestamp 1636968456
transform 1 0 17572 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_181
timestamp 1636968456
transform 1 0 18676 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_193
timestamp 1636968456
transform 1 0 19780 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_205
timestamp 1636968456
transform 1 0 20884 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_217
timestamp 1
transform 1 0 21988 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_223
timestamp 1
transform 1 0 22540 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_225
timestamp 1636968456
transform 1 0 22724 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_237
timestamp 1636968456
transform 1 0 23828 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_249
timestamp 1636968456
transform 1 0 24932 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_261
timestamp 1636968456
transform 1 0 26036 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_273
timestamp 1
transform 1 0 27140 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_279
timestamp 1
transform 1 0 27692 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_281
timestamp 1636968456
transform 1 0 27876 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_293
timestamp 1636968456
transform 1 0 28980 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_305
timestamp 1636968456
transform 1 0 30084 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_317
timestamp 1636968456
transform 1 0 31188 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_329
timestamp 1
transform 1 0 32292 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_335
timestamp 1
transform 1 0 32844 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_337
timestamp 1636968456
transform 1 0 33028 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_349
timestamp 1636968456
transform 1 0 34132 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_361
timestamp 1636968456
transform 1 0 35236 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_373
timestamp 1636968456
transform 1 0 36340 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_385
timestamp 1
transform 1 0 37444 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_391
timestamp 1
transform 1 0 37996 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_393
timestamp 1636968456
transform 1 0 38180 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_405
timestamp 1636968456
transform 1 0 39284 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_417
timestamp 1636968456
transform 1 0 40388 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_429
timestamp 1636968456
transform 1 0 41492 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_441
timestamp 1
transform 1 0 42596 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_447
timestamp 1
transform 1 0 43148 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_449
timestamp 1636968456
transform 1 0 43332 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_461
timestamp 1636968456
transform 1 0 44436 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_473
timestamp 1636968456
transform 1 0 45540 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_485
timestamp 1636968456
transform 1 0 46644 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_497
timestamp 1
transform 1 0 47748 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_503
timestamp 1
transform 1 0 48300 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_505
timestamp 1636968456
transform 1 0 48484 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_517
timestamp 1636968456
transform 1 0 49588 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_529
timestamp 1636968456
transform 1 0 50692 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_541
timestamp 1636968456
transform 1 0 51796 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_553
timestamp 1
transform 1 0 52900 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_559
timestamp 1
transform 1 0 53452 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_561
timestamp 1636968456
transform 1 0 53636 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_573
timestamp 1636968456
transform 1 0 54740 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_585
timestamp 1636968456
transform 1 0 55844 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_597
timestamp 1636968456
transform 1 0 56948 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_609
timestamp 1
transform 1 0 58052 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_615
timestamp 1
transform 1 0 58604 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_617
timestamp 1636968456
transform 1 0 58788 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_629
timestamp 1636968456
transform 1 0 59892 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_641
timestamp 1636968456
transform 1 0 60996 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_653
timestamp 1636968456
transform 1 0 62100 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_665
timestamp 1
transform 1 0 63204 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_671
timestamp 1
transform 1 0 63756 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_673
timestamp 1636968456
transform 1 0 63940 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_685
timestamp 1636968456
transform 1 0 65044 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_697
timestamp 1636968456
transform 1 0 66148 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_709
timestamp 1636968456
transform 1 0 67252 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_721
timestamp 1
transform 1 0 68356 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_727
timestamp 1
transform 1 0 68908 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_729
timestamp 1636968456
transform 1 0 69092 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_741
timestamp 1636968456
transform 1 0 70196 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_753
timestamp 1636968456
transform 1 0 71300 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_765
timestamp 1636968456
transform 1 0 72404 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_777
timestamp 1
transform 1 0 73508 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_783
timestamp 1
transform 1 0 74060 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_785
timestamp 1636968456
transform 1 0 74244 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_797
timestamp 1636968456
transform 1 0 75348 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_809
timestamp 1636968456
transform 1 0 76452 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_137_821
timestamp 1
transform 1 0 77556 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1636968456
transform 1 0 2300 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1636968456
transform 1 0 3404 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 1
transform 1 0 4508 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_29
timestamp 1636968456
transform 1 0 4692 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_41
timestamp 1636968456
transform 1 0 5796 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_53
timestamp 1
transform 1 0 6900 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_57
timestamp 1636968456
transform 1 0 7268 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_69
timestamp 1636968456
transform 1 0 8372 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1
transform 1 0 9476 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_85
timestamp 1636968456
transform 1 0 9844 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_97
timestamp 1636968456
transform 1 0 10948 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_109
timestamp 1
transform 1 0 12052 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_113
timestamp 1636968456
transform 1 0 12420 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_125
timestamp 1636968456
transform 1 0 13524 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_137
timestamp 1
transform 1 0 14628 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_141
timestamp 1636968456
transform 1 0 14996 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_153
timestamp 1636968456
transform 1 0 16100 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_165
timestamp 1
transform 1 0 17204 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_169
timestamp 1636968456
transform 1 0 17572 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_181
timestamp 1636968456
transform 1 0 18676 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_193
timestamp 1
transform 1 0 19780 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_197
timestamp 1636968456
transform 1 0 20148 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_209
timestamp 1636968456
transform 1 0 21252 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_221
timestamp 1
transform 1 0 22356 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_225
timestamp 1636968456
transform 1 0 22724 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_237
timestamp 1
transform 1 0 23828 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_241
timestamp 1
transform 1 0 24196 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_249
timestamp 1
transform 1 0 24932 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_253
timestamp 1636968456
transform 1 0 25300 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_265
timestamp 1636968456
transform 1 0 26404 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_277
timestamp 1
transform 1 0 27508 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_281
timestamp 1636968456
transform 1 0 27876 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_293
timestamp 1636968456
transform 1 0 28980 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_305
timestamp 1
transform 1 0 30084 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_309
timestamp 1636968456
transform 1 0 30452 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_321
timestamp 1636968456
transform 1 0 31556 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_333
timestamp 1
transform 1 0 32660 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_340
timestamp 1636968456
transform 1 0 33304 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_352
timestamp 1636968456
transform 1 0 34408 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_365
timestamp 1636968456
transform 1 0 35604 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_377
timestamp 1636968456
transform 1 0 36708 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_389
timestamp 1
transform 1 0 37812 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_393
timestamp 1636968456
transform 1 0 38180 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_405
timestamp 1
transform 1 0 39284 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_138_416
timestamp 1
transform 1 0 40296 0 1 77248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_138_421
timestamp 1636968456
transform 1 0 40756 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_433
timestamp 1
transform 1 0 41860 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_437
timestamp 1
transform 1 0 42228 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_445
timestamp 1
transform 1 0 42964 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_449
timestamp 1636968456
transform 1 0 43332 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_461
timestamp 1636968456
transform 1 0 44436 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_473
timestamp 1
transform 1 0 45540 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_477
timestamp 1636968456
transform 1 0 45908 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_489
timestamp 1636968456
transform 1 0 47012 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_501
timestamp 1
transform 1 0 48116 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_505
timestamp 1636968456
transform 1 0 48484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_517
timestamp 1
transform 1 0 49588 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_138_521
timestamp 1
transform 1 0 49956 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_138_529
timestamp 1
transform 1 0 50692 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_533
timestamp 1636968456
transform 1 0 51060 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_545
timestamp 1636968456
transform 1 0 52164 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_557
timestamp 1
transform 1 0 53268 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_138_561
timestamp 1
transform 1 0 53636 0 1 77248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_138_570
timestamp 1636968456
transform 1 0 54464 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_582
timestamp 1
transform 1 0 55568 0 1 77248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_138_589
timestamp 1636968456
transform 1 0 56212 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_601
timestamp 1636968456
transform 1 0 57316 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_613
timestamp 1
transform 1 0 58420 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_620
timestamp 1636968456
transform 1 0 59064 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_632
timestamp 1636968456
transform 1 0 60168 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_645
timestamp 1636968456
transform 1 0 61364 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_657
timestamp 1636968456
transform 1 0 62468 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_669
timestamp 1
transform 1 0 63572 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_673
timestamp 1636968456
transform 1 0 63940 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_685
timestamp 1636968456
transform 1 0 65044 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_697
timestamp 1
transform 1 0 66148 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_701
timestamp 1636968456
transform 1 0 66516 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_713
timestamp 1636968456
transform 1 0 67620 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_725
timestamp 1
transform 1 0 68724 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_729
timestamp 1636968456
transform 1 0 69092 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_741
timestamp 1636968456
transform 1 0 70196 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_753
timestamp 1
transform 1 0 71300 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_757
timestamp 1636968456
transform 1 0 71668 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_769
timestamp 1636968456
transform 1 0 72772 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_781
timestamp 1
transform 1 0 73876 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_785
timestamp 1636968456
transform 1 0 74244 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_797
timestamp 1636968456
transform 1 0 75348 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_809
timestamp 1
transform 1 0 76452 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_138_813
timestamp 1
transform 1 0 76820 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_138_821
timestamp 1
transform 1 0 77556 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 60260 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 75992 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 67252 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 58144 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 67068 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 67252 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 75072 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 62744 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform 1 0 70104 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1
transform -1 0 77648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 1
transform 1 0 77280 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1
transform 1 0 77280 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1
transform 1 0 77280 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1
transform 1 0 77280 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_139
timestamp 1
transform 1 0 2024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 77924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_140
timestamp 1
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 77924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_141
timestamp 1
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 77924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_142
timestamp 1
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 77924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_143
timestamp 1
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 77924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_144
timestamp 1
transform 1 0 2024 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 77924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_145
timestamp 1
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 77924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_146
timestamp 1
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 77924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_147
timestamp 1
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 77924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_148
timestamp 1
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 77924 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_149
timestamp 1
transform 1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 77924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_150
timestamp 1
transform 1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 77924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_151
timestamp 1
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 77924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_152
timestamp 1
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 77924 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_153
timestamp 1
transform 1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 77924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_154
timestamp 1
transform 1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 77924 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_155
timestamp 1
transform 1 0 2024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 77924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_156
timestamp 1
transform 1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 77924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_157
timestamp 1
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 77924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_158
timestamp 1
transform 1 0 2024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 77924 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_159
timestamp 1
transform 1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 77924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_160
timestamp 1
transform 1 0 2024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 77924 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_161
timestamp 1
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 77924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_162
timestamp 1
transform 1 0 2024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 77924 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_163
timestamp 1
transform 1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 77924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_164
timestamp 1
transform 1 0 2024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 77924 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_165
timestamp 1
transform 1 0 2024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 77924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_166
timestamp 1
transform 1 0 2024 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 77924 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_167
timestamp 1
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 77924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_168
timestamp 1
transform 1 0 2024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 77924 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_169
timestamp 1
transform 1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 77924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_170
timestamp 1
transform 1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 77924 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_171
timestamp 1
transform 1 0 2024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 77924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_172
timestamp 1
transform 1 0 2024 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 77924 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_173
timestamp 1
transform 1 0 2024 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 77924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_174
timestamp 1
transform 1 0 2024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 77924 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_175
timestamp 1
transform 1 0 2024 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 77924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_176
timestamp 1
transform 1 0 2024 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 77924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_177
timestamp 1
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 77924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_178
timestamp 1
transform 1 0 2024 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 77924 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_179
timestamp 1
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 77924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_180
timestamp 1
transform 1 0 2024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 77924 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_181
timestamp 1
transform 1 0 2024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 77924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_182
timestamp 1
transform 1 0 2024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 77924 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_183
timestamp 1
transform 1 0 2024 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 77924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_184
timestamp 1
transform 1 0 2024 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 77924 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_185
timestamp 1
transform 1 0 2024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 77924 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_186
timestamp 1
transform 1 0 2024 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 77924 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_187
timestamp 1
transform 1 0 2024 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 77924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_188
timestamp 1
transform 1 0 2024 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1
transform -1 0 77924 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_189
timestamp 1
transform 1 0 2024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1
transform -1 0 77924 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_190
timestamp 1
transform 1 0 2024 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1
transform -1 0 77924 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_191
timestamp 1
transform 1 0 2024 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1
transform -1 0 77924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_192
timestamp 1
transform 1 0 2024 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1
transform -1 0 77924 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_193
timestamp 1
transform 1 0 2024 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1
transform -1 0 77924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_194
timestamp 1
transform 1 0 2024 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1
transform -1 0 77924 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_195
timestamp 1
transform 1 0 2024 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1
transform -1 0 77924 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_196
timestamp 1
transform 1 0 2024 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1
transform -1 0 77924 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_197
timestamp 1
transform 1 0 2024 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1
transform -1 0 77924 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_198
timestamp 1
transform 1 0 2024 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1
transform -1 0 77924 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_199
timestamp 1
transform 1 0 2024 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1
transform -1 0 77924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_200
timestamp 1
transform 1 0 2024 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1
transform -1 0 77924 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_201
timestamp 1
transform 1 0 2024 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1
transform -1 0 77924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_202
timestamp 1
transform 1 0 2024 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1
transform -1 0 77924 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_203
timestamp 1
transform 1 0 2024 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1
transform -1 0 77924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_204
timestamp 1
transform 1 0 2024 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 1
transform -1 0 77924 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_205
timestamp 1
transform 1 0 2024 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 1
transform -1 0 77924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_206
timestamp 1
transform 1 0 2024 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 1
transform -1 0 77924 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_207
timestamp 1
transform 1 0 2024 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 1
transform -1 0 77924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_208
timestamp 1
transform 1 0 2024 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 1
transform -1 0 77924 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_209
timestamp 1
transform 1 0 2024 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 1
transform -1 0 77924 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_210
timestamp 1
transform 1 0 2024 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 1
transform -1 0 77924 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_211
timestamp 1
transform 1 0 2024 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 1
transform -1 0 77924 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_212
timestamp 1
transform 1 0 2024 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 1
transform -1 0 77924 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_213
timestamp 1
transform 1 0 2024 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 1
transform -1 0 77924 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_214
timestamp 1
transform 1 0 2024 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 1
transform -1 0 77924 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_215
timestamp 1
transform 1 0 2024 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 1
transform -1 0 77924 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_216
timestamp 1
transform 1 0 2024 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 1
transform -1 0 77924 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Left_217
timestamp 1
transform 1 0 2024 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_Right_78
timestamp 1
transform -1 0 77924 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Left_218
timestamp 1
transform 1 0 2024 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_Right_79
timestamp 1
transform -1 0 77924 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Left_219
timestamp 1
transform 1 0 2024 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_Right_80
timestamp 1
transform -1 0 77924 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Left_220
timestamp 1
transform 1 0 2024 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_Right_81
timestamp 1
transform -1 0 77924 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Left_221
timestamp 1
transform 1 0 2024 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_Right_82
timestamp 1
transform -1 0 77924 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Left_222
timestamp 1
transform 1 0 2024 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_Right_83
timestamp 1
transform -1 0 77924 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Left_223
timestamp 1
transform 1 0 2024 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_Right_84
timestamp 1
transform -1 0 77924 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Left_224
timestamp 1
transform 1 0 2024 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_Right_85
timestamp 1
transform -1 0 77924 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Left_225
timestamp 1
transform 1 0 2024 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_Right_86
timestamp 1
transform -1 0 77924 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Left_226
timestamp 1
transform 1 0 2024 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_Right_87
timestamp 1
transform -1 0 77924 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Left_227
timestamp 1
transform 1 0 2024 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_Right_88
timestamp 1
transform -1 0 77924 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Left_228
timestamp 1
transform 1 0 2024 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_Right_89
timestamp 1
transform -1 0 77924 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Left_229
timestamp 1
transform 1 0 2024 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_Right_90
timestamp 1
transform -1 0 77924 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Left_230
timestamp 1
transform 1 0 2024 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_Right_91
timestamp 1
transform -1 0 77924 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Left_231
timestamp 1
transform 1 0 2024 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_Right_92
timestamp 1
transform -1 0 77924 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Left_232
timestamp 1
transform 1 0 2024 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_Right_93
timestamp 1
transform -1 0 77924 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Left_233
timestamp 1
transform 1 0 2024 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_Right_94
timestamp 1
transform -1 0 77924 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Left_234
timestamp 1
transform 1 0 2024 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_Right_95
timestamp 1
transform -1 0 77924 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Left_235
timestamp 1
transform 1 0 2024 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_Right_96
timestamp 1
transform -1 0 77924 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Left_236
timestamp 1
transform 1 0 2024 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_Right_97
timestamp 1
transform -1 0 77924 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Left_237
timestamp 1
transform 1 0 2024 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_Right_98
timestamp 1
transform -1 0 77924 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Left_238
timestamp 1
transform 1 0 2024 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_Right_99
timestamp 1
transform -1 0 77924 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Left_239
timestamp 1
transform 1 0 2024 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_Right_100
timestamp 1
transform -1 0 77924 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Left_240
timestamp 1
transform 1 0 2024 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_Right_101
timestamp 1
transform -1 0 77924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_Left_241
timestamp 1
transform 1 0 2024 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_Right_102
timestamp 1
transform -1 0 77924 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_Left_242
timestamp 1
transform 1 0 2024 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_Right_103
timestamp 1
transform -1 0 77924 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_Left_243
timestamp 1
transform 1 0 2024 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_Right_104
timestamp 1
transform -1 0 77924 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_Left_244
timestamp 1
transform 1 0 2024 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_Right_105
timestamp 1
transform -1 0 77924 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Left_245
timestamp 1
transform 1 0 2024 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Right_106
timestamp 1
transform -1 0 77924 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Left_246
timestamp 1
transform 1 0 2024 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Right_107
timestamp 1
transform -1 0 77924 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Left_247
timestamp 1
transform 1 0 2024 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Right_108
timestamp 1
transform -1 0 77924 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Left_248
timestamp 1
transform 1 0 2024 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Right_109
timestamp 1
transform -1 0 77924 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Left_249
timestamp 1
transform 1 0 2024 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Right_110
timestamp 1
transform -1 0 77924 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Left_250
timestamp 1
transform 1 0 2024 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Right_111
timestamp 1
transform -1 0 77924 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Left_251
timestamp 1
transform 1 0 2024 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Right_112
timestamp 1
transform -1 0 77924 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Left_252
timestamp 1
transform 1 0 2024 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Right_113
timestamp 1
transform -1 0 77924 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Left_253
timestamp 1
transform 1 0 2024 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Right_114
timestamp 1
transform -1 0 77924 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Left_254
timestamp 1
transform 1 0 2024 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Right_115
timestamp 1
transform -1 0 77924 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Left_255
timestamp 1
transform 1 0 2024 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Right_116
timestamp 1
transform -1 0 77924 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Left_256
timestamp 1
transform 1 0 2024 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Right_117
timestamp 1
transform -1 0 77924 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Left_257
timestamp 1
transform 1 0 2024 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Right_118
timestamp 1
transform -1 0 77924 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Left_258
timestamp 1
transform 1 0 2024 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Right_119
timestamp 1
transform -1 0 77924 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Left_259
timestamp 1
transform 1 0 2024 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Right_120
timestamp 1
transform -1 0 77924 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Left_260
timestamp 1
transform 1 0 2024 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Right_121
timestamp 1
transform -1 0 77924 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Left_261
timestamp 1
transform 1 0 2024 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Right_122
timestamp 1
transform -1 0 77924 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Left_262
timestamp 1
transform 1 0 2024 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Right_123
timestamp 1
transform -1 0 77924 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Left_263
timestamp 1
transform 1 0 2024 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Right_124
timestamp 1
transform -1 0 77924 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Left_264
timestamp 1
transform 1 0 2024 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Right_125
timestamp 1
transform -1 0 77924 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Left_265
timestamp 1
transform 1 0 2024 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Right_126
timestamp 1
transform -1 0 77924 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Left_266
timestamp 1
transform 1 0 2024 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Right_127
timestamp 1
transform -1 0 77924 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Left_267
timestamp 1
transform 1 0 2024 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Right_128
timestamp 1
transform -1 0 77924 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Left_268
timestamp 1
transform 1 0 2024 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Right_129
timestamp 1
transform -1 0 77924 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Left_269
timestamp 1
transform 1 0 2024 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Right_130
timestamp 1
transform -1 0 77924 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_Left_270
timestamp 1
transform 1 0 2024 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_Right_131
timestamp 1
transform -1 0 77924 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_Left_271
timestamp 1
transform 1 0 2024 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_Right_132
timestamp 1
transform -1 0 77924 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_Left_272
timestamp 1
transform 1 0 2024 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_Right_133
timestamp 1
transform -1 0 77924 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_Left_273
timestamp 1
transform 1 0 2024 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_Right_134
timestamp 1
transform -1 0 77924 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_Left_274
timestamp 1
transform 1 0 2024 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_Right_135
timestamp 1
transform -1 0 77924 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_Left_275
timestamp 1
transform 1 0 2024 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_Right_136
timestamp 1
transform -1 0 77924 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_Left_276
timestamp 1
transform 1 0 2024 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_Right_137
timestamp 1
transform -1 0 77924 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_Left_277
timestamp 1
transform 1 0 2024 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_Right_138
timestamp 1
transform -1 0 77924 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_278
timestamp 1
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_279
timestamp 1
transform 1 0 7176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_280
timestamp 1
transform 1 0 9752 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_281
timestamp 1
transform 1 0 12328 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_282
timestamp 1
transform 1 0 14904 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_283
timestamp 1
transform 1 0 17480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_284
timestamp 1
transform 1 0 20056 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_285
timestamp 1
transform 1 0 22632 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_286
timestamp 1
transform 1 0 25208 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_287
timestamp 1
transform 1 0 27784 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_288
timestamp 1
transform 1 0 30360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_289
timestamp 1
transform 1 0 32936 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_290
timestamp 1
transform 1 0 35512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_291
timestamp 1
transform 1 0 38088 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_292
timestamp 1
transform 1 0 40664 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_293
timestamp 1
transform 1 0 43240 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_294
timestamp 1
transform 1 0 45816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_295
timestamp 1
transform 1 0 48392 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_296
timestamp 1
transform 1 0 50968 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_297
timestamp 1
transform 1 0 53544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_298
timestamp 1
transform 1 0 56120 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_299
timestamp 1
transform 1 0 58696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_300
timestamp 1
transform 1 0 61272 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_301
timestamp 1
transform 1 0 63848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_302
timestamp 1
transform 1 0 66424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_303
timestamp 1
transform 1 0 69000 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_304
timestamp 1
transform 1 0 71576 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_305
timestamp 1
transform 1 0 74152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_306
timestamp 1
transform 1 0 76728 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_307
timestamp 1
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_308
timestamp 1
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_309
timestamp 1
transform 1 0 17480 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_310
timestamp 1
transform 1 0 22632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_311
timestamp 1
transform 1 0 27784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_312
timestamp 1
transform 1 0 32936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_313
timestamp 1
transform 1 0 38088 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_314
timestamp 1
transform 1 0 43240 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_315
timestamp 1
transform 1 0 48392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_316
timestamp 1
transform 1 0 53544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_317
timestamp 1
transform 1 0 58696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_318
timestamp 1
transform 1 0 63848 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_319
timestamp 1
transform 1 0 69000 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_320
timestamp 1
transform 1 0 74152 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_321
timestamp 1
transform 1 0 4600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_322
timestamp 1
transform 1 0 9752 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_323
timestamp 1
transform 1 0 14904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_324
timestamp 1
transform 1 0 20056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_325
timestamp 1
transform 1 0 25208 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_326
timestamp 1
transform 1 0 30360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_327
timestamp 1
transform 1 0 35512 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_328
timestamp 1
transform 1 0 40664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_329
timestamp 1
transform 1 0 45816 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_330
timestamp 1
transform 1 0 50968 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_331
timestamp 1
transform 1 0 56120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_332
timestamp 1
transform 1 0 61272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_333
timestamp 1
transform 1 0 66424 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_334
timestamp 1
transform 1 0 71576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_335
timestamp 1
transform 1 0 76728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_336
timestamp 1
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_337
timestamp 1
transform 1 0 12328 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_338
timestamp 1
transform 1 0 17480 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_339
timestamp 1
transform 1 0 22632 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_340
timestamp 1
transform 1 0 27784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_341
timestamp 1
transform 1 0 32936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_342
timestamp 1
transform 1 0 38088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_343
timestamp 1
transform 1 0 43240 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_344
timestamp 1
transform 1 0 48392 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_345
timestamp 1
transform 1 0 53544 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_346
timestamp 1
transform 1 0 58696 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_347
timestamp 1
transform 1 0 63848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_348
timestamp 1
transform 1 0 69000 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_349
timestamp 1
transform 1 0 74152 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_350
timestamp 1
transform 1 0 4600 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_351
timestamp 1
transform 1 0 9752 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_352
timestamp 1
transform 1 0 14904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_353
timestamp 1
transform 1 0 20056 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_354
timestamp 1
transform 1 0 25208 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_355
timestamp 1
transform 1 0 30360 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_356
timestamp 1
transform 1 0 35512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_357
timestamp 1
transform 1 0 40664 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_358
timestamp 1
transform 1 0 45816 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_359
timestamp 1
transform 1 0 50968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_360
timestamp 1
transform 1 0 56120 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_361
timestamp 1
transform 1 0 61272 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_362
timestamp 1
transform 1 0 66424 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_363
timestamp 1
transform 1 0 71576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_364
timestamp 1
transform 1 0 76728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_365
timestamp 1
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_366
timestamp 1
transform 1 0 12328 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_367
timestamp 1
transform 1 0 17480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_368
timestamp 1
transform 1 0 22632 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_369
timestamp 1
transform 1 0 27784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_370
timestamp 1
transform 1 0 32936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_371
timestamp 1
transform 1 0 38088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_372
timestamp 1
transform 1 0 43240 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_373
timestamp 1
transform 1 0 48392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_374
timestamp 1
transform 1 0 53544 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_375
timestamp 1
transform 1 0 58696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_376
timestamp 1
transform 1 0 63848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_377
timestamp 1
transform 1 0 69000 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_378
timestamp 1
transform 1 0 74152 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_379
timestamp 1
transform 1 0 4600 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_380
timestamp 1
transform 1 0 9752 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_381
timestamp 1
transform 1 0 14904 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_382
timestamp 1
transform 1 0 20056 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_383
timestamp 1
transform 1 0 25208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_384
timestamp 1
transform 1 0 30360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_385
timestamp 1
transform 1 0 35512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_386
timestamp 1
transform 1 0 40664 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_387
timestamp 1
transform 1 0 45816 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_388
timestamp 1
transform 1 0 50968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_389
timestamp 1
transform 1 0 56120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_390
timestamp 1
transform 1 0 61272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_391
timestamp 1
transform 1 0 66424 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_392
timestamp 1
transform 1 0 71576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_393
timestamp 1
transform 1 0 76728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_394
timestamp 1
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_395
timestamp 1
transform 1 0 12328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_396
timestamp 1
transform 1 0 17480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_397
timestamp 1
transform 1 0 22632 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_398
timestamp 1
transform 1 0 27784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_399
timestamp 1
transform 1 0 32936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_400
timestamp 1
transform 1 0 38088 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_401
timestamp 1
transform 1 0 43240 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_402
timestamp 1
transform 1 0 48392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_403
timestamp 1
transform 1 0 53544 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_404
timestamp 1
transform 1 0 58696 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_405
timestamp 1
transform 1 0 63848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_406
timestamp 1
transform 1 0 69000 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_407
timestamp 1
transform 1 0 74152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_408
timestamp 1
transform 1 0 4600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_409
timestamp 1
transform 1 0 9752 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_410
timestamp 1
transform 1 0 14904 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_411
timestamp 1
transform 1 0 20056 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_412
timestamp 1
transform 1 0 25208 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_413
timestamp 1
transform 1 0 30360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_414
timestamp 1
transform 1 0 35512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_415
timestamp 1
transform 1 0 40664 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_416
timestamp 1
transform 1 0 45816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_417
timestamp 1
transform 1 0 50968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_418
timestamp 1
transform 1 0 56120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_419
timestamp 1
transform 1 0 61272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_420
timestamp 1
transform 1 0 66424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_421
timestamp 1
transform 1 0 71576 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_422
timestamp 1
transform 1 0 76728 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_423
timestamp 1
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_424
timestamp 1
transform 1 0 12328 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_425
timestamp 1
transform 1 0 17480 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_426
timestamp 1
transform 1 0 22632 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_427
timestamp 1
transform 1 0 27784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_428
timestamp 1
transform 1 0 32936 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_429
timestamp 1
transform 1 0 38088 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_430
timestamp 1
transform 1 0 43240 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_431
timestamp 1
transform 1 0 48392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_432
timestamp 1
transform 1 0 53544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_433
timestamp 1
transform 1 0 58696 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_434
timestamp 1
transform 1 0 63848 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_435
timestamp 1
transform 1 0 69000 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_436
timestamp 1
transform 1 0 74152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_437
timestamp 1
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_438
timestamp 1
transform 1 0 9752 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_439
timestamp 1
transform 1 0 14904 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_440
timestamp 1
transform 1 0 20056 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_441
timestamp 1
transform 1 0 25208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_442
timestamp 1
transform 1 0 30360 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_443
timestamp 1
transform 1 0 35512 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_444
timestamp 1
transform 1 0 40664 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_445
timestamp 1
transform 1 0 45816 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_446
timestamp 1
transform 1 0 50968 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_447
timestamp 1
transform 1 0 56120 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_448
timestamp 1
transform 1 0 61272 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_449
timestamp 1
transform 1 0 66424 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_450
timestamp 1
transform 1 0 71576 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_451
timestamp 1
transform 1 0 76728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_452
timestamp 1
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_453
timestamp 1
transform 1 0 12328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_454
timestamp 1
transform 1 0 17480 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_455
timestamp 1
transform 1 0 22632 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_456
timestamp 1
transform 1 0 27784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_457
timestamp 1
transform 1 0 32936 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_458
timestamp 1
transform 1 0 38088 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_459
timestamp 1
transform 1 0 43240 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_460
timestamp 1
transform 1 0 48392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_461
timestamp 1
transform 1 0 53544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_462
timestamp 1
transform 1 0 58696 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_463
timestamp 1
transform 1 0 63848 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_464
timestamp 1
transform 1 0 69000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_465
timestamp 1
transform 1 0 74152 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_466
timestamp 1
transform 1 0 4600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_467
timestamp 1
transform 1 0 9752 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_468
timestamp 1
transform 1 0 14904 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_469
timestamp 1
transform 1 0 20056 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_470
timestamp 1
transform 1 0 25208 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_471
timestamp 1
transform 1 0 30360 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_472
timestamp 1
transform 1 0 35512 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_473
timestamp 1
transform 1 0 40664 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_474
timestamp 1
transform 1 0 45816 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_475
timestamp 1
transform 1 0 50968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_476
timestamp 1
transform 1 0 56120 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_477
timestamp 1
transform 1 0 61272 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_478
timestamp 1
transform 1 0 66424 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_479
timestamp 1
transform 1 0 71576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_480
timestamp 1
transform 1 0 76728 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_481
timestamp 1
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_482
timestamp 1
transform 1 0 12328 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_483
timestamp 1
transform 1 0 17480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_484
timestamp 1
transform 1 0 22632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_485
timestamp 1
transform 1 0 27784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_486
timestamp 1
transform 1 0 32936 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_487
timestamp 1
transform 1 0 38088 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_488
timestamp 1
transform 1 0 43240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_489
timestamp 1
transform 1 0 48392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_490
timestamp 1
transform 1 0 53544 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_491
timestamp 1
transform 1 0 58696 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_492
timestamp 1
transform 1 0 63848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_493
timestamp 1
transform 1 0 69000 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_494
timestamp 1
transform 1 0 74152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_495
timestamp 1
transform 1 0 4600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_496
timestamp 1
transform 1 0 9752 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_497
timestamp 1
transform 1 0 14904 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_498
timestamp 1
transform 1 0 20056 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_499
timestamp 1
transform 1 0 25208 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_500
timestamp 1
transform 1 0 30360 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_501
timestamp 1
transform 1 0 35512 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_502
timestamp 1
transform 1 0 40664 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_503
timestamp 1
transform 1 0 45816 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_504
timestamp 1
transform 1 0 50968 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_505
timestamp 1
transform 1 0 56120 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_506
timestamp 1
transform 1 0 61272 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_507
timestamp 1
transform 1 0 66424 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_508
timestamp 1
transform 1 0 71576 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_509
timestamp 1
transform 1 0 76728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_510
timestamp 1
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_511
timestamp 1
transform 1 0 12328 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_512
timestamp 1
transform 1 0 17480 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_513
timestamp 1
transform 1 0 22632 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_514
timestamp 1
transform 1 0 27784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_515
timestamp 1
transform 1 0 32936 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_516
timestamp 1
transform 1 0 38088 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_517
timestamp 1
transform 1 0 43240 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_518
timestamp 1
transform 1 0 48392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_519
timestamp 1
transform 1 0 53544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_520
timestamp 1
transform 1 0 58696 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_521
timestamp 1
transform 1 0 63848 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_522
timestamp 1
transform 1 0 69000 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_523
timestamp 1
transform 1 0 74152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_524
timestamp 1
transform 1 0 4600 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_525
timestamp 1
transform 1 0 9752 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_526
timestamp 1
transform 1 0 14904 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_527
timestamp 1
transform 1 0 20056 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_528
timestamp 1
transform 1 0 25208 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_529
timestamp 1
transform 1 0 30360 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_530
timestamp 1
transform 1 0 35512 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_531
timestamp 1
transform 1 0 40664 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_532
timestamp 1
transform 1 0 45816 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_533
timestamp 1
transform 1 0 50968 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_534
timestamp 1
transform 1 0 56120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_535
timestamp 1
transform 1 0 61272 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_536
timestamp 1
transform 1 0 66424 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_537
timestamp 1
transform 1 0 71576 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_538
timestamp 1
transform 1 0 76728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_539
timestamp 1
transform 1 0 7176 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_540
timestamp 1
transform 1 0 12328 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_541
timestamp 1
transform 1 0 17480 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_542
timestamp 1
transform 1 0 22632 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_543
timestamp 1
transform 1 0 27784 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_544
timestamp 1
transform 1 0 32936 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_545
timestamp 1
transform 1 0 38088 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_546
timestamp 1
transform 1 0 43240 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_547
timestamp 1
transform 1 0 48392 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_548
timestamp 1
transform 1 0 53544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_549
timestamp 1
transform 1 0 58696 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_550
timestamp 1
transform 1 0 63848 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_551
timestamp 1
transform 1 0 69000 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_552
timestamp 1
transform 1 0 74152 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_553
timestamp 1
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_554
timestamp 1
transform 1 0 9752 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_555
timestamp 1
transform 1 0 14904 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_556
timestamp 1
transform 1 0 20056 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_557
timestamp 1
transform 1 0 25208 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_558
timestamp 1
transform 1 0 30360 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_559
timestamp 1
transform 1 0 35512 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_560
timestamp 1
transform 1 0 40664 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_561
timestamp 1
transform 1 0 45816 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_562
timestamp 1
transform 1 0 50968 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_563
timestamp 1
transform 1 0 56120 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_564
timestamp 1
transform 1 0 61272 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_565
timestamp 1
transform 1 0 66424 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_566
timestamp 1
transform 1 0 71576 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_567
timestamp 1
transform 1 0 76728 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_568
timestamp 1
transform 1 0 7176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_569
timestamp 1
transform 1 0 12328 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_570
timestamp 1
transform 1 0 17480 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_571
timestamp 1
transform 1 0 22632 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_572
timestamp 1
transform 1 0 27784 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_573
timestamp 1
transform 1 0 32936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_574
timestamp 1
transform 1 0 38088 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_575
timestamp 1
transform 1 0 43240 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_576
timestamp 1
transform 1 0 48392 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_577
timestamp 1
transform 1 0 53544 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_578
timestamp 1
transform 1 0 58696 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_579
timestamp 1
transform 1 0 63848 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_580
timestamp 1
transform 1 0 69000 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_581
timestamp 1
transform 1 0 74152 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_582
timestamp 1
transform 1 0 4600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_583
timestamp 1
transform 1 0 9752 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_584
timestamp 1
transform 1 0 14904 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_585
timestamp 1
transform 1 0 20056 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_586
timestamp 1
transform 1 0 25208 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_587
timestamp 1
transform 1 0 30360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_588
timestamp 1
transform 1 0 35512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_589
timestamp 1
transform 1 0 40664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_590
timestamp 1
transform 1 0 45816 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_591
timestamp 1
transform 1 0 50968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_592
timestamp 1
transform 1 0 56120 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_593
timestamp 1
transform 1 0 61272 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_594
timestamp 1
transform 1 0 66424 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_595
timestamp 1
transform 1 0 71576 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_596
timestamp 1
transform 1 0 76728 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_597
timestamp 1
transform 1 0 7176 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_598
timestamp 1
transform 1 0 12328 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_599
timestamp 1
transform 1 0 17480 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_600
timestamp 1
transform 1 0 22632 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_601
timestamp 1
transform 1 0 27784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_602
timestamp 1
transform 1 0 32936 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_603
timestamp 1
transform 1 0 38088 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_604
timestamp 1
transform 1 0 43240 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_605
timestamp 1
transform 1 0 48392 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_606
timestamp 1
transform 1 0 53544 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_607
timestamp 1
transform 1 0 58696 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_608
timestamp 1
transform 1 0 63848 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_609
timestamp 1
transform 1 0 69000 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_610
timestamp 1
transform 1 0 74152 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_611
timestamp 1
transform 1 0 4600 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_612
timestamp 1
transform 1 0 9752 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_613
timestamp 1
transform 1 0 14904 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_614
timestamp 1
transform 1 0 20056 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_615
timestamp 1
transform 1 0 25208 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_616
timestamp 1
transform 1 0 30360 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_617
timestamp 1
transform 1 0 35512 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_618
timestamp 1
transform 1 0 40664 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_619
timestamp 1
transform 1 0 45816 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_620
timestamp 1
transform 1 0 50968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_621
timestamp 1
transform 1 0 56120 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_622
timestamp 1
transform 1 0 61272 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_623
timestamp 1
transform 1 0 66424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_624
timestamp 1
transform 1 0 71576 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_625
timestamp 1
transform 1 0 76728 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_626
timestamp 1
transform 1 0 7176 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_627
timestamp 1
transform 1 0 12328 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_628
timestamp 1
transform 1 0 17480 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_629
timestamp 1
transform 1 0 22632 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_630
timestamp 1
transform 1 0 27784 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_631
timestamp 1
transform 1 0 32936 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_632
timestamp 1
transform 1 0 38088 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_633
timestamp 1
transform 1 0 43240 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_634
timestamp 1
transform 1 0 48392 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_635
timestamp 1
transform 1 0 53544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_636
timestamp 1
transform 1 0 58696 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_637
timestamp 1
transform 1 0 63848 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_638
timestamp 1
transform 1 0 69000 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_639
timestamp 1
transform 1 0 74152 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_640
timestamp 1
transform 1 0 4600 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_641
timestamp 1
transform 1 0 9752 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_642
timestamp 1
transform 1 0 14904 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_643
timestamp 1
transform 1 0 20056 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_644
timestamp 1
transform 1 0 25208 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_645
timestamp 1
transform 1 0 30360 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_646
timestamp 1
transform 1 0 35512 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_647
timestamp 1
transform 1 0 40664 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_648
timestamp 1
transform 1 0 45816 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_649
timestamp 1
transform 1 0 50968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_650
timestamp 1
transform 1 0 56120 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_651
timestamp 1
transform 1 0 61272 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_652
timestamp 1
transform 1 0 66424 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_653
timestamp 1
transform 1 0 71576 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_654
timestamp 1
transform 1 0 76728 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_655
timestamp 1
transform 1 0 7176 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_656
timestamp 1
transform 1 0 12328 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_657
timestamp 1
transform 1 0 17480 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_658
timestamp 1
transform 1 0 22632 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_659
timestamp 1
transform 1 0 27784 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_660
timestamp 1
transform 1 0 32936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_661
timestamp 1
transform 1 0 38088 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_662
timestamp 1
transform 1 0 43240 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_663
timestamp 1
transform 1 0 48392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_664
timestamp 1
transform 1 0 53544 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_665
timestamp 1
transform 1 0 58696 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_666
timestamp 1
transform 1 0 63848 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_667
timestamp 1
transform 1 0 69000 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_668
timestamp 1
transform 1 0 74152 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_669
timestamp 1
transform 1 0 4600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_670
timestamp 1
transform 1 0 9752 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_671
timestamp 1
transform 1 0 14904 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_672
timestamp 1
transform 1 0 20056 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_673
timestamp 1
transform 1 0 25208 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_674
timestamp 1
transform 1 0 30360 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_675
timestamp 1
transform 1 0 35512 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_676
timestamp 1
transform 1 0 40664 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_677
timestamp 1
transform 1 0 45816 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_678
timestamp 1
transform 1 0 50968 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_679
timestamp 1
transform 1 0 56120 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_680
timestamp 1
transform 1 0 61272 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_681
timestamp 1
transform 1 0 66424 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_682
timestamp 1
transform 1 0 71576 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_683
timestamp 1
transform 1 0 76728 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_684
timestamp 1
transform 1 0 7176 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_685
timestamp 1
transform 1 0 12328 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_686
timestamp 1
transform 1 0 17480 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_687
timestamp 1
transform 1 0 22632 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_688
timestamp 1
transform 1 0 27784 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_689
timestamp 1
transform 1 0 32936 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_690
timestamp 1
transform 1 0 38088 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_691
timestamp 1
transform 1 0 43240 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_692
timestamp 1
transform 1 0 48392 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_693
timestamp 1
transform 1 0 53544 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_694
timestamp 1
transform 1 0 58696 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_695
timestamp 1
transform 1 0 63848 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_696
timestamp 1
transform 1 0 69000 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_697
timestamp 1
transform 1 0 74152 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_698
timestamp 1
transform 1 0 4600 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_699
timestamp 1
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_700
timestamp 1
transform 1 0 14904 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_701
timestamp 1
transform 1 0 20056 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_702
timestamp 1
transform 1 0 25208 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_703
timestamp 1
transform 1 0 30360 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_704
timestamp 1
transform 1 0 35512 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_705
timestamp 1
transform 1 0 40664 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_706
timestamp 1
transform 1 0 45816 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_707
timestamp 1
transform 1 0 50968 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_708
timestamp 1
transform 1 0 56120 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_709
timestamp 1
transform 1 0 61272 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_710
timestamp 1
transform 1 0 66424 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_711
timestamp 1
transform 1 0 71576 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_712
timestamp 1
transform 1 0 76728 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_713
timestamp 1
transform 1 0 7176 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_714
timestamp 1
transform 1 0 12328 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_715
timestamp 1
transform 1 0 17480 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_716
timestamp 1
transform 1 0 22632 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_717
timestamp 1
transform 1 0 27784 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_718
timestamp 1
transform 1 0 32936 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_719
timestamp 1
transform 1 0 38088 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_720
timestamp 1
transform 1 0 43240 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_721
timestamp 1
transform 1 0 48392 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_722
timestamp 1
transform 1 0 53544 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_723
timestamp 1
transform 1 0 58696 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_724
timestamp 1
transform 1 0 63848 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_725
timestamp 1
transform 1 0 69000 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_726
timestamp 1
transform 1 0 74152 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_727
timestamp 1
transform 1 0 4600 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_728
timestamp 1
transform 1 0 9752 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_729
timestamp 1
transform 1 0 14904 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_730
timestamp 1
transform 1 0 20056 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_731
timestamp 1
transform 1 0 25208 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_732
timestamp 1
transform 1 0 30360 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_733
timestamp 1
transform 1 0 35512 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_734
timestamp 1
transform 1 0 40664 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_735
timestamp 1
transform 1 0 45816 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_736
timestamp 1
transform 1 0 50968 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_737
timestamp 1
transform 1 0 56120 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_738
timestamp 1
transform 1 0 61272 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_739
timestamp 1
transform 1 0 66424 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_740
timestamp 1
transform 1 0 71576 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_741
timestamp 1
transform 1 0 76728 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_742
timestamp 1
transform 1 0 7176 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_743
timestamp 1
transform 1 0 12328 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_744
timestamp 1
transform 1 0 17480 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_745
timestamp 1
transform 1 0 22632 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_746
timestamp 1
transform 1 0 27784 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_747
timestamp 1
transform 1 0 32936 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_748
timestamp 1
transform 1 0 38088 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_749
timestamp 1
transform 1 0 43240 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_750
timestamp 1
transform 1 0 48392 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_751
timestamp 1
transform 1 0 53544 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_752
timestamp 1
transform 1 0 58696 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_753
timestamp 1
transform 1 0 63848 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_754
timestamp 1
transform 1 0 69000 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_755
timestamp 1
transform 1 0 74152 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_756
timestamp 1
transform 1 0 4600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_757
timestamp 1
transform 1 0 9752 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_758
timestamp 1
transform 1 0 14904 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_759
timestamp 1
transform 1 0 20056 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_760
timestamp 1
transform 1 0 25208 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_761
timestamp 1
transform 1 0 30360 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_762
timestamp 1
transform 1 0 35512 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_763
timestamp 1
transform 1 0 40664 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_764
timestamp 1
transform 1 0 45816 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_765
timestamp 1
transform 1 0 50968 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_766
timestamp 1
transform 1 0 56120 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_767
timestamp 1
transform 1 0 61272 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_768
timestamp 1
transform 1 0 66424 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_769
timestamp 1
transform 1 0 71576 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_770
timestamp 1
transform 1 0 76728 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_771
timestamp 1
transform 1 0 7176 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_772
timestamp 1
transform 1 0 12328 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_773
timestamp 1
transform 1 0 17480 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_774
timestamp 1
transform 1 0 22632 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_775
timestamp 1
transform 1 0 27784 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_776
timestamp 1
transform 1 0 32936 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_777
timestamp 1
transform 1 0 38088 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_778
timestamp 1
transform 1 0 43240 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_779
timestamp 1
transform 1 0 48392 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_780
timestamp 1
transform 1 0 53544 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_781
timestamp 1
transform 1 0 58696 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_782
timestamp 1
transform 1 0 63848 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_783
timestamp 1
transform 1 0 69000 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_784
timestamp 1
transform 1 0 74152 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_785
timestamp 1
transform 1 0 4600 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_786
timestamp 1
transform 1 0 9752 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_787
timestamp 1
transform 1 0 14904 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_788
timestamp 1
transform 1 0 20056 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_789
timestamp 1
transform 1 0 25208 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_790
timestamp 1
transform 1 0 30360 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_791
timestamp 1
transform 1 0 35512 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_792
timestamp 1
transform 1 0 40664 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_793
timestamp 1
transform 1 0 45816 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_794
timestamp 1
transform 1 0 50968 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_795
timestamp 1
transform 1 0 56120 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_796
timestamp 1
transform 1 0 61272 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_797
timestamp 1
transform 1 0 66424 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_798
timestamp 1
transform 1 0 71576 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_799
timestamp 1
transform 1 0 76728 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_800
timestamp 1
transform 1 0 7176 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_801
timestamp 1
transform 1 0 12328 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_802
timestamp 1
transform 1 0 17480 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_803
timestamp 1
transform 1 0 22632 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_804
timestamp 1
transform 1 0 27784 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_805
timestamp 1
transform 1 0 32936 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_806
timestamp 1
transform 1 0 38088 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_807
timestamp 1
transform 1 0 43240 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_808
timestamp 1
transform 1 0 48392 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_809
timestamp 1
transform 1 0 53544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_810
timestamp 1
transform 1 0 58696 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_811
timestamp 1
transform 1 0 63848 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_812
timestamp 1
transform 1 0 69000 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_813
timestamp 1
transform 1 0 74152 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_814
timestamp 1
transform 1 0 4600 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_815
timestamp 1
transform 1 0 9752 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_816
timestamp 1
transform 1 0 14904 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_817
timestamp 1
transform 1 0 20056 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_818
timestamp 1
transform 1 0 25208 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_819
timestamp 1
transform 1 0 30360 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_820
timestamp 1
transform 1 0 35512 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_821
timestamp 1
transform 1 0 40664 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_822
timestamp 1
transform 1 0 45816 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_823
timestamp 1
transform 1 0 50968 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_824
timestamp 1
transform 1 0 56120 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_825
timestamp 1
transform 1 0 61272 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_826
timestamp 1
transform 1 0 66424 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_827
timestamp 1
transform 1 0 71576 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_828
timestamp 1
transform 1 0 76728 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_829
timestamp 1
transform 1 0 7176 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_830
timestamp 1
transform 1 0 12328 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_831
timestamp 1
transform 1 0 17480 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_832
timestamp 1
transform 1 0 22632 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_833
timestamp 1
transform 1 0 27784 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_834
timestamp 1
transform 1 0 32936 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_835
timestamp 1
transform 1 0 38088 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_836
timestamp 1
transform 1 0 43240 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_837
timestamp 1
transform 1 0 48392 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_838
timestamp 1
transform 1 0 53544 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_839
timestamp 1
transform 1 0 58696 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_840
timestamp 1
transform 1 0 63848 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_841
timestamp 1
transform 1 0 69000 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_842
timestamp 1
transform 1 0 74152 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_843
timestamp 1
transform 1 0 4600 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_844
timestamp 1
transform 1 0 9752 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_845
timestamp 1
transform 1 0 14904 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_846
timestamp 1
transform 1 0 20056 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_847
timestamp 1
transform 1 0 25208 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_848
timestamp 1
transform 1 0 30360 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_849
timestamp 1
transform 1 0 35512 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_850
timestamp 1
transform 1 0 40664 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_851
timestamp 1
transform 1 0 45816 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_852
timestamp 1
transform 1 0 50968 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_853
timestamp 1
transform 1 0 56120 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_854
timestamp 1
transform 1 0 61272 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_855
timestamp 1
transform 1 0 66424 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_856
timestamp 1
transform 1 0 71576 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_857
timestamp 1
transform 1 0 76728 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_858
timestamp 1
transform 1 0 7176 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_859
timestamp 1
transform 1 0 12328 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_860
timestamp 1
transform 1 0 17480 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_861
timestamp 1
transform 1 0 22632 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_862
timestamp 1
transform 1 0 27784 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_863
timestamp 1
transform 1 0 32936 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_864
timestamp 1
transform 1 0 38088 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_865
timestamp 1
transform 1 0 43240 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_866
timestamp 1
transform 1 0 48392 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_867
timestamp 1
transform 1 0 53544 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_868
timestamp 1
transform 1 0 58696 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_869
timestamp 1
transform 1 0 63848 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_870
timestamp 1
transform 1 0 69000 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_871
timestamp 1
transform 1 0 74152 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_872
timestamp 1
transform 1 0 4600 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_873
timestamp 1
transform 1 0 9752 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_874
timestamp 1
transform 1 0 14904 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_875
timestamp 1
transform 1 0 20056 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_876
timestamp 1
transform 1 0 25208 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_877
timestamp 1
transform 1 0 30360 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_878
timestamp 1
transform 1 0 35512 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_879
timestamp 1
transform 1 0 40664 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_880
timestamp 1
transform 1 0 45816 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_881
timestamp 1
transform 1 0 50968 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_882
timestamp 1
transform 1 0 56120 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_883
timestamp 1
transform 1 0 61272 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_884
timestamp 1
transform 1 0 66424 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_885
timestamp 1
transform 1 0 71576 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_886
timestamp 1
transform 1 0 76728 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_887
timestamp 1
transform 1 0 7176 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_888
timestamp 1
transform 1 0 12328 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_889
timestamp 1
transform 1 0 17480 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_890
timestamp 1
transform 1 0 22632 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_891
timestamp 1
transform 1 0 27784 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_892
timestamp 1
transform 1 0 32936 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_893
timestamp 1
transform 1 0 38088 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_894
timestamp 1
transform 1 0 43240 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_895
timestamp 1
transform 1 0 48392 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_896
timestamp 1
transform 1 0 53544 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_897
timestamp 1
transform 1 0 58696 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_898
timestamp 1
transform 1 0 63848 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_899
timestamp 1
transform 1 0 69000 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_900
timestamp 1
transform 1 0 74152 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_901
timestamp 1
transform 1 0 4600 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_902
timestamp 1
transform 1 0 9752 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_903
timestamp 1
transform 1 0 14904 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_904
timestamp 1
transform 1 0 20056 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_905
timestamp 1
transform 1 0 25208 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_906
timestamp 1
transform 1 0 30360 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_907
timestamp 1
transform 1 0 35512 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_908
timestamp 1
transform 1 0 40664 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_909
timestamp 1
transform 1 0 45816 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_910
timestamp 1
transform 1 0 50968 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_911
timestamp 1
transform 1 0 56120 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_912
timestamp 1
transform 1 0 61272 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_913
timestamp 1
transform 1 0 66424 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_914
timestamp 1
transform 1 0 71576 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_915
timestamp 1
transform 1 0 76728 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_916
timestamp 1
transform 1 0 7176 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_917
timestamp 1
transform 1 0 12328 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_918
timestamp 1
transform 1 0 17480 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_919
timestamp 1
transform 1 0 22632 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_920
timestamp 1
transform 1 0 27784 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_921
timestamp 1
transform 1 0 32936 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_922
timestamp 1
transform 1 0 38088 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_923
timestamp 1
transform 1 0 43240 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_924
timestamp 1
transform 1 0 48392 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_925
timestamp 1
transform 1 0 53544 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_926
timestamp 1
transform 1 0 58696 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_927
timestamp 1
transform 1 0 63848 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_928
timestamp 1
transform 1 0 69000 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_929
timestamp 1
transform 1 0 74152 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_930
timestamp 1
transform 1 0 4600 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_931
timestamp 1
transform 1 0 9752 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_932
timestamp 1
transform 1 0 14904 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_933
timestamp 1
transform 1 0 20056 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_934
timestamp 1
transform 1 0 25208 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_935
timestamp 1
transform 1 0 30360 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_936
timestamp 1
transform 1 0 35512 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_937
timestamp 1
transform 1 0 40664 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_938
timestamp 1
transform 1 0 45816 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_939
timestamp 1
transform 1 0 50968 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_940
timestamp 1
transform 1 0 56120 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_941
timestamp 1
transform 1 0 61272 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_942
timestamp 1
transform 1 0 66424 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_943
timestamp 1
transform 1 0 71576 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_944
timestamp 1
transform 1 0 76728 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_945
timestamp 1
transform 1 0 7176 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_946
timestamp 1
transform 1 0 12328 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_947
timestamp 1
transform 1 0 17480 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_948
timestamp 1
transform 1 0 22632 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_949
timestamp 1
transform 1 0 27784 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_950
timestamp 1
transform 1 0 32936 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_951
timestamp 1
transform 1 0 38088 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_952
timestamp 1
transform 1 0 43240 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_953
timestamp 1
transform 1 0 48392 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_954
timestamp 1
transform 1 0 53544 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_955
timestamp 1
transform 1 0 58696 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_956
timestamp 1
transform 1 0 63848 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_957
timestamp 1
transform 1 0 69000 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_958
timestamp 1
transform 1 0 74152 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_959
timestamp 1
transform 1 0 4600 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_960
timestamp 1
transform 1 0 9752 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_961
timestamp 1
transform 1 0 14904 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_962
timestamp 1
transform 1 0 20056 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_963
timestamp 1
transform 1 0 25208 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_964
timestamp 1
transform 1 0 30360 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_965
timestamp 1
transform 1 0 35512 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_966
timestamp 1
transform 1 0 40664 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_967
timestamp 1
transform 1 0 45816 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_968
timestamp 1
transform 1 0 50968 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_969
timestamp 1
transform 1 0 56120 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_970
timestamp 1
transform 1 0 61272 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_971
timestamp 1
transform 1 0 66424 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_972
timestamp 1
transform 1 0 71576 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_973
timestamp 1
transform 1 0 76728 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_974
timestamp 1
transform 1 0 7176 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_975
timestamp 1
transform 1 0 12328 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_976
timestamp 1
transform 1 0 17480 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_977
timestamp 1
transform 1 0 22632 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_978
timestamp 1
transform 1 0 27784 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_979
timestamp 1
transform 1 0 32936 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_980
timestamp 1
transform 1 0 38088 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_981
timestamp 1
transform 1 0 43240 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_982
timestamp 1
transform 1 0 48392 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_983
timestamp 1
transform 1 0 53544 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_984
timestamp 1
transform 1 0 58696 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_985
timestamp 1
transform 1 0 63848 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_986
timestamp 1
transform 1 0 69000 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_987
timestamp 1
transform 1 0 74152 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_988
timestamp 1
transform 1 0 4600 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_989
timestamp 1
transform 1 0 9752 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_990
timestamp 1
transform 1 0 14904 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_991
timestamp 1
transform 1 0 20056 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_992
timestamp 1
transform 1 0 25208 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_993
timestamp 1
transform 1 0 30360 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_994
timestamp 1
transform 1 0 35512 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_995
timestamp 1
transform 1 0 40664 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_996
timestamp 1
transform 1 0 45816 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_997
timestamp 1
transform 1 0 50968 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_998
timestamp 1
transform 1 0 56120 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_999
timestamp 1
transform 1 0 61272 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1000
timestamp 1
transform 1 0 66424 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1001
timestamp 1
transform 1 0 71576 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1002
timestamp 1
transform 1 0 76728 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1003
timestamp 1
transform 1 0 7176 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1004
timestamp 1
transform 1 0 12328 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1005
timestamp 1
transform 1 0 17480 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1006
timestamp 1
transform 1 0 22632 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1007
timestamp 1
transform 1 0 27784 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1008
timestamp 1
transform 1 0 32936 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1009
timestamp 1
transform 1 0 38088 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1010
timestamp 1
transform 1 0 43240 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1011
timestamp 1
transform 1 0 48392 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1012
timestamp 1
transform 1 0 53544 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1013
timestamp 1
transform 1 0 58696 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1014
timestamp 1
transform 1 0 63848 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1015
timestamp 1
transform 1 0 69000 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_1016
timestamp 1
transform 1 0 74152 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1017
timestamp 1
transform 1 0 4600 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1018
timestamp 1
transform 1 0 9752 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1019
timestamp 1
transform 1 0 14904 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1020
timestamp 1
transform 1 0 20056 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1021
timestamp 1
transform 1 0 25208 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1022
timestamp 1
transform 1 0 30360 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1023
timestamp 1
transform 1 0 35512 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1024
timestamp 1
transform 1 0 40664 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1025
timestamp 1
transform 1 0 45816 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1026
timestamp 1
transform 1 0 50968 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1027
timestamp 1
transform 1 0 56120 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1028
timestamp 1
transform 1 0 61272 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1029
timestamp 1
transform 1 0 66424 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1030
timestamp 1
transform 1 0 71576 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1031
timestamp 1
transform 1 0 76728 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1032
timestamp 1
transform 1 0 7176 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1033
timestamp 1
transform 1 0 12328 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1034
timestamp 1
transform 1 0 17480 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1035
timestamp 1
transform 1 0 22632 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1036
timestamp 1
transform 1 0 27784 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1037
timestamp 1
transform 1 0 32936 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1038
timestamp 1
transform 1 0 38088 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1039
timestamp 1
transform 1 0 43240 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1040
timestamp 1
transform 1 0 48392 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1041
timestamp 1
transform 1 0 53544 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1042
timestamp 1
transform 1 0 58696 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1043
timestamp 1
transform 1 0 63848 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1044
timestamp 1
transform 1 0 69000 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_1045
timestamp 1
transform 1 0 74152 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1046
timestamp 1
transform 1 0 4600 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1047
timestamp 1
transform 1 0 9752 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1048
timestamp 1
transform 1 0 14904 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1049
timestamp 1
transform 1 0 20056 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1050
timestamp 1
transform 1 0 25208 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1051
timestamp 1
transform 1 0 30360 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1052
timestamp 1
transform 1 0 35512 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1053
timestamp 1
transform 1 0 40664 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1054
timestamp 1
transform 1 0 45816 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1055
timestamp 1
transform 1 0 50968 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1056
timestamp 1
transform 1 0 56120 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1057
timestamp 1
transform 1 0 61272 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1058
timestamp 1
transform 1 0 66424 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1059
timestamp 1
transform 1 0 71576 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1060
timestamp 1
transform 1 0 76728 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1061
timestamp 1
transform 1 0 7176 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1062
timestamp 1
transform 1 0 12328 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1063
timestamp 1
transform 1 0 17480 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1064
timestamp 1
transform 1 0 22632 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1065
timestamp 1
transform 1 0 27784 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1066
timestamp 1
transform 1 0 32936 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1067
timestamp 1
transform 1 0 38088 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1068
timestamp 1
transform 1 0 43240 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1069
timestamp 1
transform 1 0 48392 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1070
timestamp 1
transform 1 0 53544 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1071
timestamp 1
transform 1 0 58696 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1072
timestamp 1
transform 1 0 63848 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1073
timestamp 1
transform 1 0 69000 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_1074
timestamp 1
transform 1 0 74152 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1075
timestamp 1
transform 1 0 4600 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1076
timestamp 1
transform 1 0 9752 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1077
timestamp 1
transform 1 0 14904 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1078
timestamp 1
transform 1 0 20056 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1079
timestamp 1
transform 1 0 25208 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1080
timestamp 1
transform 1 0 30360 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1081
timestamp 1
transform 1 0 35512 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1082
timestamp 1
transform 1 0 40664 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1083
timestamp 1
transform 1 0 45816 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1084
timestamp 1
transform 1 0 50968 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1085
timestamp 1
transform 1 0 56120 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1086
timestamp 1
transform 1 0 61272 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1087
timestamp 1
transform 1 0 66424 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1088
timestamp 1
transform 1 0 71576 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1089
timestamp 1
transform 1 0 76728 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1090
timestamp 1
transform 1 0 7176 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1091
timestamp 1
transform 1 0 12328 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1092
timestamp 1
transform 1 0 17480 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1093
timestamp 1
transform 1 0 22632 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1094
timestamp 1
transform 1 0 27784 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1095
timestamp 1
transform 1 0 32936 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1096
timestamp 1
transform 1 0 38088 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1097
timestamp 1
transform 1 0 43240 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1098
timestamp 1
transform 1 0 48392 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1099
timestamp 1
transform 1 0 53544 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1100
timestamp 1
transform 1 0 58696 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1101
timestamp 1
transform 1 0 63848 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1102
timestamp 1
transform 1 0 69000 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_1103
timestamp 1
transform 1 0 74152 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1104
timestamp 1
transform 1 0 4600 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1105
timestamp 1
transform 1 0 9752 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1106
timestamp 1
transform 1 0 14904 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1107
timestamp 1
transform 1 0 20056 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1108
timestamp 1
transform 1 0 25208 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1109
timestamp 1
transform 1 0 30360 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1110
timestamp 1
transform 1 0 35512 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1111
timestamp 1
transform 1 0 40664 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1112
timestamp 1
transform 1 0 45816 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1113
timestamp 1
transform 1 0 50968 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1114
timestamp 1
transform 1 0 56120 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1115
timestamp 1
transform 1 0 61272 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1116
timestamp 1
transform 1 0 66424 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1117
timestamp 1
transform 1 0 71576 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1118
timestamp 1
transform 1 0 76728 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1119
timestamp 1
transform 1 0 7176 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1120
timestamp 1
transform 1 0 12328 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1121
timestamp 1
transform 1 0 17480 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1122
timestamp 1
transform 1 0 22632 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1123
timestamp 1
transform 1 0 27784 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1124
timestamp 1
transform 1 0 32936 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1125
timestamp 1
transform 1 0 38088 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1126
timestamp 1
transform 1 0 43240 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1127
timestamp 1
transform 1 0 48392 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1128
timestamp 1
transform 1 0 53544 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1129
timestamp 1
transform 1 0 58696 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1130
timestamp 1
transform 1 0 63848 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1131
timestamp 1
transform 1 0 69000 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_1132
timestamp 1
transform 1 0 74152 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1133
timestamp 1
transform 1 0 4600 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1134
timestamp 1
transform 1 0 9752 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1135
timestamp 1
transform 1 0 14904 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1136
timestamp 1
transform 1 0 20056 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1137
timestamp 1
transform 1 0 25208 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1138
timestamp 1
transform 1 0 30360 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1139
timestamp 1
transform 1 0 35512 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1140
timestamp 1
transform 1 0 40664 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1141
timestamp 1
transform 1 0 45816 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1142
timestamp 1
transform 1 0 50968 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1143
timestamp 1
transform 1 0 56120 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1144
timestamp 1
transform 1 0 61272 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1145
timestamp 1
transform 1 0 66424 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1146
timestamp 1
transform 1 0 71576 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1147
timestamp 1
transform 1 0 76728 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1148
timestamp 1
transform 1 0 7176 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1149
timestamp 1
transform 1 0 12328 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1150
timestamp 1
transform 1 0 17480 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1151
timestamp 1
transform 1 0 22632 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1152
timestamp 1
transform 1 0 27784 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1153
timestamp 1
transform 1 0 32936 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1154
timestamp 1
transform 1 0 38088 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1155
timestamp 1
transform 1 0 43240 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1156
timestamp 1
transform 1 0 48392 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1157
timestamp 1
transform 1 0 53544 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1158
timestamp 1
transform 1 0 58696 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1159
timestamp 1
transform 1 0 63848 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1160
timestamp 1
transform 1 0 69000 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_1161
timestamp 1
transform 1 0 74152 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1162
timestamp 1
transform 1 0 4600 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1163
timestamp 1
transform 1 0 9752 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1164
timestamp 1
transform 1 0 14904 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1165
timestamp 1
transform 1 0 20056 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1166
timestamp 1
transform 1 0 25208 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1167
timestamp 1
transform 1 0 30360 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1168
timestamp 1
transform 1 0 35512 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1169
timestamp 1
transform 1 0 40664 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1170
timestamp 1
transform 1 0 45816 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1171
timestamp 1
transform 1 0 50968 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1172
timestamp 1
transform 1 0 56120 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1173
timestamp 1
transform 1 0 61272 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1174
timestamp 1
transform 1 0 66424 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1175
timestamp 1
transform 1 0 71576 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1176
timestamp 1
transform 1 0 76728 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1177
timestamp 1
transform 1 0 7176 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1178
timestamp 1
transform 1 0 12328 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1179
timestamp 1
transform 1 0 17480 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1180
timestamp 1
transform 1 0 22632 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1181
timestamp 1
transform 1 0 27784 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1182
timestamp 1
transform 1 0 32936 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1183
timestamp 1
transform 1 0 38088 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1184
timestamp 1
transform 1 0 43240 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1185
timestamp 1
transform 1 0 48392 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1186
timestamp 1
transform 1 0 53544 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1187
timestamp 1
transform 1 0 58696 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1188
timestamp 1
transform 1 0 63848 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1189
timestamp 1
transform 1 0 69000 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_1190
timestamp 1
transform 1 0 74152 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1191
timestamp 1
transform 1 0 4600 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1192
timestamp 1
transform 1 0 9752 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1193
timestamp 1
transform 1 0 14904 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1194
timestamp 1
transform 1 0 20056 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1195
timestamp 1
transform 1 0 25208 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1196
timestamp 1
transform 1 0 30360 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1197
timestamp 1
transform 1 0 35512 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1198
timestamp 1
transform 1 0 40664 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1199
timestamp 1
transform 1 0 45816 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1200
timestamp 1
transform 1 0 50968 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1201
timestamp 1
transform 1 0 56120 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1202
timestamp 1
transform 1 0 61272 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1203
timestamp 1
transform 1 0 66424 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1204
timestamp 1
transform 1 0 71576 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1205
timestamp 1
transform 1 0 76728 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1206
timestamp 1
transform 1 0 7176 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1207
timestamp 1
transform 1 0 12328 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1208
timestamp 1
transform 1 0 17480 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1209
timestamp 1
transform 1 0 22632 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1210
timestamp 1
transform 1 0 27784 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1211
timestamp 1
transform 1 0 32936 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1212
timestamp 1
transform 1 0 38088 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1213
timestamp 1
transform 1 0 43240 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1214
timestamp 1
transform 1 0 48392 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1215
timestamp 1
transform 1 0 53544 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1216
timestamp 1
transform 1 0 58696 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1217
timestamp 1
transform 1 0 63848 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1218
timestamp 1
transform 1 0 69000 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_1219
timestamp 1
transform 1 0 74152 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1220
timestamp 1
transform 1 0 4600 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1221
timestamp 1
transform 1 0 9752 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1222
timestamp 1
transform 1 0 14904 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1223
timestamp 1
transform 1 0 20056 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1224
timestamp 1
transform 1 0 25208 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1225
timestamp 1
transform 1 0 30360 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1226
timestamp 1
transform 1 0 35512 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1227
timestamp 1
transform 1 0 40664 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1228
timestamp 1
transform 1 0 45816 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1229
timestamp 1
transform 1 0 50968 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1230
timestamp 1
transform 1 0 56120 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1231
timestamp 1
transform 1 0 61272 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1232
timestamp 1
transform 1 0 66424 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1233
timestamp 1
transform 1 0 71576 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1234
timestamp 1
transform 1 0 76728 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1235
timestamp 1
transform 1 0 7176 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1236
timestamp 1
transform 1 0 12328 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1237
timestamp 1
transform 1 0 17480 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1238
timestamp 1
transform 1 0 22632 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1239
timestamp 1
transform 1 0 27784 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1240
timestamp 1
transform 1 0 32936 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1241
timestamp 1
transform 1 0 38088 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1242
timestamp 1
transform 1 0 43240 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1243
timestamp 1
transform 1 0 48392 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1244
timestamp 1
transform 1 0 53544 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1245
timestamp 1
transform 1 0 58696 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1246
timestamp 1
transform 1 0 63848 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1247
timestamp 1
transform 1 0 69000 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_1248
timestamp 1
transform 1 0 74152 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1249
timestamp 1
transform 1 0 4600 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1250
timestamp 1
transform 1 0 9752 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1251
timestamp 1
transform 1 0 14904 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1252
timestamp 1
transform 1 0 20056 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1253
timestamp 1
transform 1 0 25208 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1254
timestamp 1
transform 1 0 30360 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1255
timestamp 1
transform 1 0 35512 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1256
timestamp 1
transform 1 0 40664 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1257
timestamp 1
transform 1 0 45816 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1258
timestamp 1
transform 1 0 50968 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1259
timestamp 1
transform 1 0 56120 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1260
timestamp 1
transform 1 0 61272 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1261
timestamp 1
transform 1 0 66424 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1262
timestamp 1
transform 1 0 71576 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1263
timestamp 1
transform 1 0 76728 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1264
timestamp 1
transform 1 0 7176 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1265
timestamp 1
transform 1 0 12328 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1266
timestamp 1
transform 1 0 17480 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1267
timestamp 1
transform 1 0 22632 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1268
timestamp 1
transform 1 0 27784 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1269
timestamp 1
transform 1 0 32936 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1270
timestamp 1
transform 1 0 38088 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1271
timestamp 1
transform 1 0 43240 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1272
timestamp 1
transform 1 0 48392 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1273
timestamp 1
transform 1 0 53544 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1274
timestamp 1
transform 1 0 58696 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1275
timestamp 1
transform 1 0 63848 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1276
timestamp 1
transform 1 0 69000 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_1277
timestamp 1
transform 1 0 74152 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1278
timestamp 1
transform 1 0 4600 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1279
timestamp 1
transform 1 0 9752 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1280
timestamp 1
transform 1 0 14904 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1281
timestamp 1
transform 1 0 20056 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1282
timestamp 1
transform 1 0 25208 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1283
timestamp 1
transform 1 0 30360 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1284
timestamp 1
transform 1 0 35512 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1285
timestamp 1
transform 1 0 40664 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1286
timestamp 1
transform 1 0 45816 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1287
timestamp 1
transform 1 0 50968 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1288
timestamp 1
transform 1 0 56120 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1289
timestamp 1
transform 1 0 61272 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1290
timestamp 1
transform 1 0 66424 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1291
timestamp 1
transform 1 0 71576 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1292
timestamp 1
transform 1 0 76728 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1293
timestamp 1
transform 1 0 7176 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1294
timestamp 1
transform 1 0 12328 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1295
timestamp 1
transform 1 0 17480 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1296
timestamp 1
transform 1 0 22632 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1297
timestamp 1
transform 1 0 27784 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1298
timestamp 1
transform 1 0 32936 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1299
timestamp 1
transform 1 0 38088 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1300
timestamp 1
transform 1 0 43240 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1301
timestamp 1
transform 1 0 48392 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1302
timestamp 1
transform 1 0 53544 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1303
timestamp 1
transform 1 0 58696 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1304
timestamp 1
transform 1 0 63848 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1305
timestamp 1
transform 1 0 69000 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_1306
timestamp 1
transform 1 0 74152 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1307
timestamp 1
transform 1 0 4600 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1308
timestamp 1
transform 1 0 9752 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1309
timestamp 1
transform 1 0 14904 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1310
timestamp 1
transform 1 0 20056 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1311
timestamp 1
transform 1 0 25208 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1312
timestamp 1
transform 1 0 30360 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1313
timestamp 1
transform 1 0 35512 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1314
timestamp 1
transform 1 0 40664 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1315
timestamp 1
transform 1 0 45816 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1316
timestamp 1
transform 1 0 50968 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1317
timestamp 1
transform 1 0 56120 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1318
timestamp 1
transform 1 0 61272 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1319
timestamp 1
transform 1 0 66424 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1320
timestamp 1
transform 1 0 71576 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1321
timestamp 1
transform 1 0 76728 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1322
timestamp 1
transform 1 0 7176 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1323
timestamp 1
transform 1 0 12328 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1324
timestamp 1
transform 1 0 17480 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1325
timestamp 1
transform 1 0 22632 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1326
timestamp 1
transform 1 0 27784 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1327
timestamp 1
transform 1 0 32936 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1328
timestamp 1
transform 1 0 38088 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1329
timestamp 1
transform 1 0 43240 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1330
timestamp 1
transform 1 0 48392 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1331
timestamp 1
transform 1 0 53544 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1332
timestamp 1
transform 1 0 58696 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1333
timestamp 1
transform 1 0 63848 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1334
timestamp 1
transform 1 0 69000 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_1335
timestamp 1
transform 1 0 74152 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1336
timestamp 1
transform 1 0 4600 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1337
timestamp 1
transform 1 0 9752 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1338
timestamp 1
transform 1 0 14904 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1339
timestamp 1
transform 1 0 20056 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1340
timestamp 1
transform 1 0 25208 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1341
timestamp 1
transform 1 0 30360 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1342
timestamp 1
transform 1 0 35512 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1343
timestamp 1
transform 1 0 40664 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1344
timestamp 1
transform 1 0 45816 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1345
timestamp 1
transform 1 0 50968 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1346
timestamp 1
transform 1 0 56120 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1347
timestamp 1
transform 1 0 61272 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1348
timestamp 1
transform 1 0 66424 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1349
timestamp 1
transform 1 0 71576 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1350
timestamp 1
transform 1 0 76728 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1351
timestamp 1
transform 1 0 7176 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1352
timestamp 1
transform 1 0 12328 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1353
timestamp 1
transform 1 0 17480 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1354
timestamp 1
transform 1 0 22632 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1355
timestamp 1
transform 1 0 27784 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1356
timestamp 1
transform 1 0 32936 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1357
timestamp 1
transform 1 0 38088 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1358
timestamp 1
transform 1 0 43240 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1359
timestamp 1
transform 1 0 48392 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1360
timestamp 1
transform 1 0 53544 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1361
timestamp 1
transform 1 0 58696 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1362
timestamp 1
transform 1 0 63848 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1363
timestamp 1
transform 1 0 69000 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_1364
timestamp 1
transform 1 0 74152 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1365
timestamp 1
transform 1 0 4600 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1366
timestamp 1
transform 1 0 9752 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1367
timestamp 1
transform 1 0 14904 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1368
timestamp 1
transform 1 0 20056 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1369
timestamp 1
transform 1 0 25208 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1370
timestamp 1
transform 1 0 30360 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1371
timestamp 1
transform 1 0 35512 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1372
timestamp 1
transform 1 0 40664 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1373
timestamp 1
transform 1 0 45816 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1374
timestamp 1
transform 1 0 50968 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1375
timestamp 1
transform 1 0 56120 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1376
timestamp 1
transform 1 0 61272 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1377
timestamp 1
transform 1 0 66424 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1378
timestamp 1
transform 1 0 71576 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1379
timestamp 1
transform 1 0 76728 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1380
timestamp 1
transform 1 0 7176 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1381
timestamp 1
transform 1 0 12328 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1382
timestamp 1
transform 1 0 17480 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1383
timestamp 1
transform 1 0 22632 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1384
timestamp 1
transform 1 0 27784 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1385
timestamp 1
transform 1 0 32936 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1386
timestamp 1
transform 1 0 38088 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1387
timestamp 1
transform 1 0 43240 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1388
timestamp 1
transform 1 0 48392 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1389
timestamp 1
transform 1 0 53544 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1390
timestamp 1
transform 1 0 58696 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1391
timestamp 1
transform 1 0 63848 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1392
timestamp 1
transform 1 0 69000 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_1393
timestamp 1
transform 1 0 74152 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1394
timestamp 1
transform 1 0 4600 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1395
timestamp 1
transform 1 0 9752 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1396
timestamp 1
transform 1 0 14904 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1397
timestamp 1
transform 1 0 20056 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1398
timestamp 1
transform 1 0 25208 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1399
timestamp 1
transform 1 0 30360 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1400
timestamp 1
transform 1 0 35512 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1401
timestamp 1
transform 1 0 40664 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1402
timestamp 1
transform 1 0 45816 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1403
timestamp 1
transform 1 0 50968 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1404
timestamp 1
transform 1 0 56120 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1405
timestamp 1
transform 1 0 61272 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1406
timestamp 1
transform 1 0 66424 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1407
timestamp 1
transform 1 0 71576 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1408
timestamp 1
transform 1 0 76728 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1409
timestamp 1
transform 1 0 7176 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1410
timestamp 1
transform 1 0 12328 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1411
timestamp 1
transform 1 0 17480 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1412
timestamp 1
transform 1 0 22632 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1413
timestamp 1
transform 1 0 27784 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1414
timestamp 1
transform 1 0 32936 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1415
timestamp 1
transform 1 0 38088 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1416
timestamp 1
transform 1 0 43240 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1417
timestamp 1
transform 1 0 48392 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1418
timestamp 1
transform 1 0 53544 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1419
timestamp 1
transform 1 0 58696 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1420
timestamp 1
transform 1 0 63848 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1421
timestamp 1
transform 1 0 69000 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_1422
timestamp 1
transform 1 0 74152 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1423
timestamp 1
transform 1 0 4600 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1424
timestamp 1
transform 1 0 9752 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1425
timestamp 1
transform 1 0 14904 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1426
timestamp 1
transform 1 0 20056 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1427
timestamp 1
transform 1 0 25208 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1428
timestamp 1
transform 1 0 30360 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1429
timestamp 1
transform 1 0 35512 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1430
timestamp 1
transform 1 0 40664 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1431
timestamp 1
transform 1 0 45816 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1432
timestamp 1
transform 1 0 50968 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1433
timestamp 1
transform 1 0 56120 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1434
timestamp 1
transform 1 0 61272 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1435
timestamp 1
transform 1 0 66424 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1436
timestamp 1
transform 1 0 71576 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1437
timestamp 1
transform 1 0 76728 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1438
timestamp 1
transform 1 0 7176 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1439
timestamp 1
transform 1 0 12328 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1440
timestamp 1
transform 1 0 17480 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1441
timestamp 1
transform 1 0 22632 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1442
timestamp 1
transform 1 0 27784 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1443
timestamp 1
transform 1 0 32936 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1444
timestamp 1
transform 1 0 38088 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1445
timestamp 1
transform 1 0 43240 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1446
timestamp 1
transform 1 0 48392 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1447
timestamp 1
transform 1 0 53544 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1448
timestamp 1
transform 1 0 58696 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1449
timestamp 1
transform 1 0 63848 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1450
timestamp 1
transform 1 0 69000 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_79_1451
timestamp 1
transform 1 0 74152 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1452
timestamp 1
transform 1 0 4600 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1453
timestamp 1
transform 1 0 9752 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1454
timestamp 1
transform 1 0 14904 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1455
timestamp 1
transform 1 0 20056 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1456
timestamp 1
transform 1 0 25208 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1457
timestamp 1
transform 1 0 30360 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1458
timestamp 1
transform 1 0 35512 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1459
timestamp 1
transform 1 0 40664 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1460
timestamp 1
transform 1 0 45816 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1461
timestamp 1
transform 1 0 50968 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1462
timestamp 1
transform 1 0 56120 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1463
timestamp 1
transform 1 0 61272 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1464
timestamp 1
transform 1 0 66424 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1465
timestamp 1
transform 1 0 71576 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1466
timestamp 1
transform 1 0 76728 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1467
timestamp 1
transform 1 0 7176 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1468
timestamp 1
transform 1 0 12328 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1469
timestamp 1
transform 1 0 17480 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1470
timestamp 1
transform 1 0 22632 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1471
timestamp 1
transform 1 0 27784 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1472
timestamp 1
transform 1 0 32936 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1473
timestamp 1
transform 1 0 38088 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1474
timestamp 1
transform 1 0 43240 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1475
timestamp 1
transform 1 0 48392 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1476
timestamp 1
transform 1 0 53544 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1477
timestamp 1
transform 1 0 58696 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1478
timestamp 1
transform 1 0 63848 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1479
timestamp 1
transform 1 0 69000 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_81_1480
timestamp 1
transform 1 0 74152 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1481
timestamp 1
transform 1 0 4600 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1482
timestamp 1
transform 1 0 9752 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1483
timestamp 1
transform 1 0 14904 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1484
timestamp 1
transform 1 0 20056 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1485
timestamp 1
transform 1 0 25208 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1486
timestamp 1
transform 1 0 30360 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1487
timestamp 1
transform 1 0 35512 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1488
timestamp 1
transform 1 0 40664 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1489
timestamp 1
transform 1 0 45816 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1490
timestamp 1
transform 1 0 50968 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1491
timestamp 1
transform 1 0 56120 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1492
timestamp 1
transform 1 0 61272 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1493
timestamp 1
transform 1 0 66424 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1494
timestamp 1
transform 1 0 71576 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1495
timestamp 1
transform 1 0 76728 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1496
timestamp 1
transform 1 0 7176 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1497
timestamp 1
transform 1 0 12328 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1498
timestamp 1
transform 1 0 17480 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1499
timestamp 1
transform 1 0 22632 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1500
timestamp 1
transform 1 0 27784 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1501
timestamp 1
transform 1 0 32936 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1502
timestamp 1
transform 1 0 38088 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1503
timestamp 1
transform 1 0 43240 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1504
timestamp 1
transform 1 0 48392 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1505
timestamp 1
transform 1 0 53544 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1506
timestamp 1
transform 1 0 58696 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1507
timestamp 1
transform 1 0 63848 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1508
timestamp 1
transform 1 0 69000 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_83_1509
timestamp 1
transform 1 0 74152 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1510
timestamp 1
transform 1 0 4600 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1511
timestamp 1
transform 1 0 9752 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1512
timestamp 1
transform 1 0 14904 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1513
timestamp 1
transform 1 0 20056 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1514
timestamp 1
transform 1 0 25208 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1515
timestamp 1
transform 1 0 30360 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1516
timestamp 1
transform 1 0 35512 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1517
timestamp 1
transform 1 0 40664 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1518
timestamp 1
transform 1 0 45816 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1519
timestamp 1
transform 1 0 50968 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1520
timestamp 1
transform 1 0 56120 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1521
timestamp 1
transform 1 0 61272 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1522
timestamp 1
transform 1 0 66424 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1523
timestamp 1
transform 1 0 71576 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1524
timestamp 1
transform 1 0 76728 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1525
timestamp 1
transform 1 0 7176 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1526
timestamp 1
transform 1 0 12328 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1527
timestamp 1
transform 1 0 17480 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1528
timestamp 1
transform 1 0 22632 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1529
timestamp 1
transform 1 0 27784 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1530
timestamp 1
transform 1 0 32936 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1531
timestamp 1
transform 1 0 38088 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1532
timestamp 1
transform 1 0 43240 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1533
timestamp 1
transform 1 0 48392 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1534
timestamp 1
transform 1 0 53544 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1535
timestamp 1
transform 1 0 58696 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1536
timestamp 1
transform 1 0 63848 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1537
timestamp 1
transform 1 0 69000 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_85_1538
timestamp 1
transform 1 0 74152 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1539
timestamp 1
transform 1 0 4600 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1540
timestamp 1
transform 1 0 9752 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1541
timestamp 1
transform 1 0 14904 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1542
timestamp 1
transform 1 0 20056 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1543
timestamp 1
transform 1 0 25208 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1544
timestamp 1
transform 1 0 30360 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1545
timestamp 1
transform 1 0 35512 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1546
timestamp 1
transform 1 0 40664 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1547
timestamp 1
transform 1 0 45816 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1548
timestamp 1
transform 1 0 50968 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1549
timestamp 1
transform 1 0 56120 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1550
timestamp 1
transform 1 0 61272 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1551
timestamp 1
transform 1 0 66424 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1552
timestamp 1
transform 1 0 71576 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1553
timestamp 1
transform 1 0 76728 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1554
timestamp 1
transform 1 0 7176 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1555
timestamp 1
transform 1 0 12328 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1556
timestamp 1
transform 1 0 17480 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1557
timestamp 1
transform 1 0 22632 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1558
timestamp 1
transform 1 0 27784 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1559
timestamp 1
transform 1 0 32936 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1560
timestamp 1
transform 1 0 38088 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1561
timestamp 1
transform 1 0 43240 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1562
timestamp 1
transform 1 0 48392 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1563
timestamp 1
transform 1 0 53544 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1564
timestamp 1
transform 1 0 58696 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1565
timestamp 1
transform 1 0 63848 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1566
timestamp 1
transform 1 0 69000 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_87_1567
timestamp 1
transform 1 0 74152 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1568
timestamp 1
transform 1 0 4600 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1569
timestamp 1
transform 1 0 9752 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1570
timestamp 1
transform 1 0 14904 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1571
timestamp 1
transform 1 0 20056 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1572
timestamp 1
transform 1 0 25208 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1573
timestamp 1
transform 1 0 30360 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1574
timestamp 1
transform 1 0 35512 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1575
timestamp 1
transform 1 0 40664 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1576
timestamp 1
transform 1 0 45816 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1577
timestamp 1
transform 1 0 50968 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1578
timestamp 1
transform 1 0 56120 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1579
timestamp 1
transform 1 0 61272 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1580
timestamp 1
transform 1 0 66424 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1581
timestamp 1
transform 1 0 71576 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1582
timestamp 1
transform 1 0 76728 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1583
timestamp 1
transform 1 0 7176 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1584
timestamp 1
transform 1 0 12328 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1585
timestamp 1
transform 1 0 17480 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1586
timestamp 1
transform 1 0 22632 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1587
timestamp 1
transform 1 0 27784 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1588
timestamp 1
transform 1 0 32936 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1589
timestamp 1
transform 1 0 38088 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1590
timestamp 1
transform 1 0 43240 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1591
timestamp 1
transform 1 0 48392 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1592
timestamp 1
transform 1 0 53544 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1593
timestamp 1
transform 1 0 58696 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1594
timestamp 1
transform 1 0 63848 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1595
timestamp 1
transform 1 0 69000 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_89_1596
timestamp 1
transform 1 0 74152 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1597
timestamp 1
transform 1 0 4600 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1598
timestamp 1
transform 1 0 9752 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1599
timestamp 1
transform 1 0 14904 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1600
timestamp 1
transform 1 0 20056 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1601
timestamp 1
transform 1 0 25208 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1602
timestamp 1
transform 1 0 30360 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1603
timestamp 1
transform 1 0 35512 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1604
timestamp 1
transform 1 0 40664 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1605
timestamp 1
transform 1 0 45816 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1606
timestamp 1
transform 1 0 50968 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1607
timestamp 1
transform 1 0 56120 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1608
timestamp 1
transform 1 0 61272 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1609
timestamp 1
transform 1 0 66424 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1610
timestamp 1
transform 1 0 71576 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1611
timestamp 1
transform 1 0 76728 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1612
timestamp 1
transform 1 0 7176 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1613
timestamp 1
transform 1 0 12328 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1614
timestamp 1
transform 1 0 17480 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1615
timestamp 1
transform 1 0 22632 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1616
timestamp 1
transform 1 0 27784 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1617
timestamp 1
transform 1 0 32936 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1618
timestamp 1
transform 1 0 38088 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1619
timestamp 1
transform 1 0 43240 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1620
timestamp 1
transform 1 0 48392 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1621
timestamp 1
transform 1 0 53544 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1622
timestamp 1
transform 1 0 58696 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1623
timestamp 1
transform 1 0 63848 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1624
timestamp 1
transform 1 0 69000 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_91_1625
timestamp 1
transform 1 0 74152 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1626
timestamp 1
transform 1 0 4600 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1627
timestamp 1
transform 1 0 9752 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1628
timestamp 1
transform 1 0 14904 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1629
timestamp 1
transform 1 0 20056 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1630
timestamp 1
transform 1 0 25208 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1631
timestamp 1
transform 1 0 30360 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1632
timestamp 1
transform 1 0 35512 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1633
timestamp 1
transform 1 0 40664 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1634
timestamp 1
transform 1 0 45816 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1635
timestamp 1
transform 1 0 50968 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1636
timestamp 1
transform 1 0 56120 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1637
timestamp 1
transform 1 0 61272 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1638
timestamp 1
transform 1 0 66424 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1639
timestamp 1
transform 1 0 71576 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1640
timestamp 1
transform 1 0 76728 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1641
timestamp 1
transform 1 0 7176 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1642
timestamp 1
transform 1 0 12328 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1643
timestamp 1
transform 1 0 17480 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1644
timestamp 1
transform 1 0 22632 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1645
timestamp 1
transform 1 0 27784 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1646
timestamp 1
transform 1 0 32936 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1647
timestamp 1
transform 1 0 38088 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1648
timestamp 1
transform 1 0 43240 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1649
timestamp 1
transform 1 0 48392 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1650
timestamp 1
transform 1 0 53544 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1651
timestamp 1
transform 1 0 58696 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1652
timestamp 1
transform 1 0 63848 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1653
timestamp 1
transform 1 0 69000 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_93_1654
timestamp 1
transform 1 0 74152 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1655
timestamp 1
transform 1 0 4600 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1656
timestamp 1
transform 1 0 9752 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1657
timestamp 1
transform 1 0 14904 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1658
timestamp 1
transform 1 0 20056 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1659
timestamp 1
transform 1 0 25208 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1660
timestamp 1
transform 1 0 30360 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1661
timestamp 1
transform 1 0 35512 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1662
timestamp 1
transform 1 0 40664 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1663
timestamp 1
transform 1 0 45816 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1664
timestamp 1
transform 1 0 50968 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1665
timestamp 1
transform 1 0 56120 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1666
timestamp 1
transform 1 0 61272 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1667
timestamp 1
transform 1 0 66424 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1668
timestamp 1
transform 1 0 71576 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1669
timestamp 1
transform 1 0 76728 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1670
timestamp 1
transform 1 0 7176 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1671
timestamp 1
transform 1 0 12328 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1672
timestamp 1
transform 1 0 17480 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1673
timestamp 1
transform 1 0 22632 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1674
timestamp 1
transform 1 0 27784 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1675
timestamp 1
transform 1 0 32936 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1676
timestamp 1
transform 1 0 38088 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1677
timestamp 1
transform 1 0 43240 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1678
timestamp 1
transform 1 0 48392 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1679
timestamp 1
transform 1 0 53544 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1680
timestamp 1
transform 1 0 58696 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1681
timestamp 1
transform 1 0 63848 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1682
timestamp 1
transform 1 0 69000 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_95_1683
timestamp 1
transform 1 0 74152 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1684
timestamp 1
transform 1 0 4600 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1685
timestamp 1
transform 1 0 9752 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1686
timestamp 1
transform 1 0 14904 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1687
timestamp 1
transform 1 0 20056 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1688
timestamp 1
transform 1 0 25208 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1689
timestamp 1
transform 1 0 30360 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1690
timestamp 1
transform 1 0 35512 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1691
timestamp 1
transform 1 0 40664 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1692
timestamp 1
transform 1 0 45816 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1693
timestamp 1
transform 1 0 50968 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1694
timestamp 1
transform 1 0 56120 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1695
timestamp 1
transform 1 0 61272 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1696
timestamp 1
transform 1 0 66424 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1697
timestamp 1
transform 1 0 71576 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1698
timestamp 1
transform 1 0 76728 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1699
timestamp 1
transform 1 0 7176 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1700
timestamp 1
transform 1 0 12328 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1701
timestamp 1
transform 1 0 17480 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1702
timestamp 1
transform 1 0 22632 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1703
timestamp 1
transform 1 0 27784 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1704
timestamp 1
transform 1 0 32936 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1705
timestamp 1
transform 1 0 38088 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1706
timestamp 1
transform 1 0 43240 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1707
timestamp 1
transform 1 0 48392 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1708
timestamp 1
transform 1 0 53544 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1709
timestamp 1
transform 1 0 58696 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1710
timestamp 1
transform 1 0 63848 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1711
timestamp 1
transform 1 0 69000 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_97_1712
timestamp 1
transform 1 0 74152 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1713
timestamp 1
transform 1 0 4600 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1714
timestamp 1
transform 1 0 9752 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1715
timestamp 1
transform 1 0 14904 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1716
timestamp 1
transform 1 0 20056 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1717
timestamp 1
transform 1 0 25208 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1718
timestamp 1
transform 1 0 30360 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1719
timestamp 1
transform 1 0 35512 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1720
timestamp 1
transform 1 0 40664 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1721
timestamp 1
transform 1 0 45816 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1722
timestamp 1
transform 1 0 50968 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1723
timestamp 1
transform 1 0 56120 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1724
timestamp 1
transform 1 0 61272 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1725
timestamp 1
transform 1 0 66424 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1726
timestamp 1
transform 1 0 71576 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1727
timestamp 1
transform 1 0 76728 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1728
timestamp 1
transform 1 0 7176 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1729
timestamp 1
transform 1 0 12328 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1730
timestamp 1
transform 1 0 17480 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1731
timestamp 1
transform 1 0 22632 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1732
timestamp 1
transform 1 0 27784 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1733
timestamp 1
transform 1 0 32936 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1734
timestamp 1
transform 1 0 38088 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1735
timestamp 1
transform 1 0 43240 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1736
timestamp 1
transform 1 0 48392 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1737
timestamp 1
transform 1 0 53544 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1738
timestamp 1
transform 1 0 58696 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1739
timestamp 1
transform 1 0 63848 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1740
timestamp 1
transform 1 0 69000 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_99_1741
timestamp 1
transform 1 0 74152 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1742
timestamp 1
transform 1 0 4600 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1743
timestamp 1
transform 1 0 9752 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1744
timestamp 1
transform 1 0 14904 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1745
timestamp 1
transform 1 0 20056 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1746
timestamp 1
transform 1 0 25208 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1747
timestamp 1
transform 1 0 30360 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1748
timestamp 1
transform 1 0 35512 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1749
timestamp 1
transform 1 0 40664 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1750
timestamp 1
transform 1 0 45816 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1751
timestamp 1
transform 1 0 50968 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1752
timestamp 1
transform 1 0 56120 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1753
timestamp 1
transform 1 0 61272 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1754
timestamp 1
transform 1 0 66424 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1755
timestamp 1
transform 1 0 71576 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1756
timestamp 1
transform 1 0 76728 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1757
timestamp 1
transform 1 0 7176 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1758
timestamp 1
transform 1 0 12328 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1759
timestamp 1
transform 1 0 17480 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1760
timestamp 1
transform 1 0 22632 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1761
timestamp 1
transform 1 0 27784 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1762
timestamp 1
transform 1 0 32936 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1763
timestamp 1
transform 1 0 38088 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1764
timestamp 1
transform 1 0 43240 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1765
timestamp 1
transform 1 0 48392 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1766
timestamp 1
transform 1 0 53544 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1767
timestamp 1
transform 1 0 58696 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1768
timestamp 1
transform 1 0 63848 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1769
timestamp 1
transform 1 0 69000 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_101_1770
timestamp 1
transform 1 0 74152 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1771
timestamp 1
transform 1 0 4600 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1772
timestamp 1
transform 1 0 9752 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1773
timestamp 1
transform 1 0 14904 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1774
timestamp 1
transform 1 0 20056 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1775
timestamp 1
transform 1 0 25208 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1776
timestamp 1
transform 1 0 30360 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1777
timestamp 1
transform 1 0 35512 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1778
timestamp 1
transform 1 0 40664 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1779
timestamp 1
transform 1 0 45816 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1780
timestamp 1
transform 1 0 50968 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1781
timestamp 1
transform 1 0 56120 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1782
timestamp 1
transform 1 0 61272 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1783
timestamp 1
transform 1 0 66424 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1784
timestamp 1
transform 1 0 71576 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1785
timestamp 1
transform 1 0 76728 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1786
timestamp 1
transform 1 0 7176 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1787
timestamp 1
transform 1 0 12328 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1788
timestamp 1
transform 1 0 17480 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1789
timestamp 1
transform 1 0 22632 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1790
timestamp 1
transform 1 0 27784 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1791
timestamp 1
transform 1 0 32936 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1792
timestamp 1
transform 1 0 38088 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1793
timestamp 1
transform 1 0 43240 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1794
timestamp 1
transform 1 0 48392 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1795
timestamp 1
transform 1 0 53544 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1796
timestamp 1
transform 1 0 58696 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1797
timestamp 1
transform 1 0 63848 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1798
timestamp 1
transform 1 0 69000 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_103_1799
timestamp 1
transform 1 0 74152 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1800
timestamp 1
transform 1 0 4600 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1801
timestamp 1
transform 1 0 9752 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1802
timestamp 1
transform 1 0 14904 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1803
timestamp 1
transform 1 0 20056 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1804
timestamp 1
transform 1 0 25208 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1805
timestamp 1
transform 1 0 30360 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1806
timestamp 1
transform 1 0 35512 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1807
timestamp 1
transform 1 0 40664 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1808
timestamp 1
transform 1 0 45816 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1809
timestamp 1
transform 1 0 50968 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1810
timestamp 1
transform 1 0 56120 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1811
timestamp 1
transform 1 0 61272 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1812
timestamp 1
transform 1 0 66424 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1813
timestamp 1
transform 1 0 71576 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1814
timestamp 1
transform 1 0 76728 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1815
timestamp 1
transform 1 0 7176 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1816
timestamp 1
transform 1 0 12328 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1817
timestamp 1
transform 1 0 17480 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1818
timestamp 1
transform 1 0 22632 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1819
timestamp 1
transform 1 0 27784 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1820
timestamp 1
transform 1 0 32936 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1821
timestamp 1
transform 1 0 38088 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1822
timestamp 1
transform 1 0 43240 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1823
timestamp 1
transform 1 0 48392 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1824
timestamp 1
transform 1 0 53544 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1825
timestamp 1
transform 1 0 58696 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1826
timestamp 1
transform 1 0 63848 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1827
timestamp 1
transform 1 0 69000 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_105_1828
timestamp 1
transform 1 0 74152 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1829
timestamp 1
transform 1 0 4600 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1830
timestamp 1
transform 1 0 9752 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1831
timestamp 1
transform 1 0 14904 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1832
timestamp 1
transform 1 0 20056 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1833
timestamp 1
transform 1 0 25208 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1834
timestamp 1
transform 1 0 30360 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1835
timestamp 1
transform 1 0 35512 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1836
timestamp 1
transform 1 0 40664 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1837
timestamp 1
transform 1 0 45816 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1838
timestamp 1
transform 1 0 50968 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1839
timestamp 1
transform 1 0 56120 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1840
timestamp 1
transform 1 0 61272 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1841
timestamp 1
transform 1 0 66424 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1842
timestamp 1
transform 1 0 71576 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1843
timestamp 1
transform 1 0 76728 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1844
timestamp 1
transform 1 0 7176 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1845
timestamp 1
transform 1 0 12328 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1846
timestamp 1
transform 1 0 17480 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1847
timestamp 1
transform 1 0 22632 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1848
timestamp 1
transform 1 0 27784 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1849
timestamp 1
transform 1 0 32936 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1850
timestamp 1
transform 1 0 38088 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1851
timestamp 1
transform 1 0 43240 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1852
timestamp 1
transform 1 0 48392 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1853
timestamp 1
transform 1 0 53544 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1854
timestamp 1
transform 1 0 58696 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1855
timestamp 1
transform 1 0 63848 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1856
timestamp 1
transform 1 0 69000 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_1857
timestamp 1
transform 1 0 74152 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1858
timestamp 1
transform 1 0 4600 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1859
timestamp 1
transform 1 0 9752 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1860
timestamp 1
transform 1 0 14904 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1861
timestamp 1
transform 1 0 20056 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1862
timestamp 1
transform 1 0 25208 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1863
timestamp 1
transform 1 0 30360 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1864
timestamp 1
transform 1 0 35512 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1865
timestamp 1
transform 1 0 40664 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1866
timestamp 1
transform 1 0 45816 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1867
timestamp 1
transform 1 0 50968 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1868
timestamp 1
transform 1 0 56120 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1869
timestamp 1
transform 1 0 61272 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1870
timestamp 1
transform 1 0 66424 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1871
timestamp 1
transform 1 0 71576 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1872
timestamp 1
transform 1 0 76728 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1873
timestamp 1
transform 1 0 7176 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1874
timestamp 1
transform 1 0 12328 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1875
timestamp 1
transform 1 0 17480 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1876
timestamp 1
transform 1 0 22632 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1877
timestamp 1
transform 1 0 27784 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1878
timestamp 1
transform 1 0 32936 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1879
timestamp 1
transform 1 0 38088 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1880
timestamp 1
transform 1 0 43240 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1881
timestamp 1
transform 1 0 48392 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1882
timestamp 1
transform 1 0 53544 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1883
timestamp 1
transform 1 0 58696 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1884
timestamp 1
transform 1 0 63848 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1885
timestamp 1
transform 1 0 69000 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_1886
timestamp 1
transform 1 0 74152 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1887
timestamp 1
transform 1 0 4600 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1888
timestamp 1
transform 1 0 9752 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1889
timestamp 1
transform 1 0 14904 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1890
timestamp 1
transform 1 0 20056 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1891
timestamp 1
transform 1 0 25208 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1892
timestamp 1
transform 1 0 30360 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1893
timestamp 1
transform 1 0 35512 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1894
timestamp 1
transform 1 0 40664 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1895
timestamp 1
transform 1 0 45816 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1896
timestamp 1
transform 1 0 50968 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1897
timestamp 1
transform 1 0 56120 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1898
timestamp 1
transform 1 0 61272 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1899
timestamp 1
transform 1 0 66424 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1900
timestamp 1
transform 1 0 71576 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1901
timestamp 1
transform 1 0 76728 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1902
timestamp 1
transform 1 0 7176 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1903
timestamp 1
transform 1 0 12328 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1904
timestamp 1
transform 1 0 17480 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1905
timestamp 1
transform 1 0 22632 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1906
timestamp 1
transform 1 0 27784 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1907
timestamp 1
transform 1 0 32936 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1908
timestamp 1
transform 1 0 38088 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1909
timestamp 1
transform 1 0 43240 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1910
timestamp 1
transform 1 0 48392 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1911
timestamp 1
transform 1 0 53544 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1912
timestamp 1
transform 1 0 58696 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1913
timestamp 1
transform 1 0 63848 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1914
timestamp 1
transform 1 0 69000 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_1915
timestamp 1
transform 1 0 74152 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1916
timestamp 1
transform 1 0 4600 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1917
timestamp 1
transform 1 0 9752 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1918
timestamp 1
transform 1 0 14904 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1919
timestamp 1
transform 1 0 20056 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1920
timestamp 1
transform 1 0 25208 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1921
timestamp 1
transform 1 0 30360 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1922
timestamp 1
transform 1 0 35512 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1923
timestamp 1
transform 1 0 40664 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1924
timestamp 1
transform 1 0 45816 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1925
timestamp 1
transform 1 0 50968 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1926
timestamp 1
transform 1 0 56120 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1927
timestamp 1
transform 1 0 61272 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1928
timestamp 1
transform 1 0 66424 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1929
timestamp 1
transform 1 0 71576 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1930
timestamp 1
transform 1 0 76728 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1931
timestamp 1
transform 1 0 7176 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1932
timestamp 1
transform 1 0 12328 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1933
timestamp 1
transform 1 0 17480 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1934
timestamp 1
transform 1 0 22632 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1935
timestamp 1
transform 1 0 27784 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1936
timestamp 1
transform 1 0 32936 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1937
timestamp 1
transform 1 0 38088 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1938
timestamp 1
transform 1 0 43240 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1939
timestamp 1
transform 1 0 48392 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1940
timestamp 1
transform 1 0 53544 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1941
timestamp 1
transform 1 0 58696 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1942
timestamp 1
transform 1 0 63848 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1943
timestamp 1
transform 1 0 69000 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_1944
timestamp 1
transform 1 0 74152 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1945
timestamp 1
transform 1 0 4600 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1946
timestamp 1
transform 1 0 9752 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1947
timestamp 1
transform 1 0 14904 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1948
timestamp 1
transform 1 0 20056 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1949
timestamp 1
transform 1 0 25208 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1950
timestamp 1
transform 1 0 30360 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1951
timestamp 1
transform 1 0 35512 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1952
timestamp 1
transform 1 0 40664 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1953
timestamp 1
transform 1 0 45816 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1954
timestamp 1
transform 1 0 50968 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1955
timestamp 1
transform 1 0 56120 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1956
timestamp 1
transform 1 0 61272 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1957
timestamp 1
transform 1 0 66424 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1958
timestamp 1
transform 1 0 71576 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1959
timestamp 1
transform 1 0 76728 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1960
timestamp 1
transform 1 0 7176 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1961
timestamp 1
transform 1 0 12328 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1962
timestamp 1
transform 1 0 17480 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1963
timestamp 1
transform 1 0 22632 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1964
timestamp 1
transform 1 0 27784 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1965
timestamp 1
transform 1 0 32936 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1966
timestamp 1
transform 1 0 38088 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1967
timestamp 1
transform 1 0 43240 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1968
timestamp 1
transform 1 0 48392 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1969
timestamp 1
transform 1 0 53544 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1970
timestamp 1
transform 1 0 58696 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1971
timestamp 1
transform 1 0 63848 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1972
timestamp 1
transform 1 0 69000 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_1973
timestamp 1
transform 1 0 74152 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1974
timestamp 1
transform 1 0 4600 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1975
timestamp 1
transform 1 0 9752 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1976
timestamp 1
transform 1 0 14904 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1977
timestamp 1
transform 1 0 20056 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1978
timestamp 1
transform 1 0 25208 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1979
timestamp 1
transform 1 0 30360 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1980
timestamp 1
transform 1 0 35512 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1981
timestamp 1
transform 1 0 40664 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1982
timestamp 1
transform 1 0 45816 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1983
timestamp 1
transform 1 0 50968 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1984
timestamp 1
transform 1 0 56120 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1985
timestamp 1
transform 1 0 61272 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1986
timestamp 1
transform 1 0 66424 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1987
timestamp 1
transform 1 0 71576 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1988
timestamp 1
transform 1 0 76728 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1989
timestamp 1
transform 1 0 7176 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1990
timestamp 1
transform 1 0 12328 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1991
timestamp 1
transform 1 0 17480 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1992
timestamp 1
transform 1 0 22632 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1993
timestamp 1
transform 1 0 27784 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1994
timestamp 1
transform 1 0 32936 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1995
timestamp 1
transform 1 0 38088 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1996
timestamp 1
transform 1 0 43240 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1997
timestamp 1
transform 1 0 48392 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1998
timestamp 1
transform 1 0 53544 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_1999
timestamp 1
transform 1 0 58696 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_2000
timestamp 1
transform 1 0 63848 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_2001
timestamp 1
transform 1 0 69000 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_2002
timestamp 1
transform 1 0 74152 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2003
timestamp 1
transform 1 0 4600 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2004
timestamp 1
transform 1 0 9752 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2005
timestamp 1
transform 1 0 14904 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2006
timestamp 1
transform 1 0 20056 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2007
timestamp 1
transform 1 0 25208 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2008
timestamp 1
transform 1 0 30360 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2009
timestamp 1
transform 1 0 35512 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2010
timestamp 1
transform 1 0 40664 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2011
timestamp 1
transform 1 0 45816 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2012
timestamp 1
transform 1 0 50968 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2013
timestamp 1
transform 1 0 56120 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2014
timestamp 1
transform 1 0 61272 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2015
timestamp 1
transform 1 0 66424 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2016
timestamp 1
transform 1 0 71576 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_2017
timestamp 1
transform 1 0 76728 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2018
timestamp 1
transform 1 0 7176 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2019
timestamp 1
transform 1 0 12328 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2020
timestamp 1
transform 1 0 17480 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2021
timestamp 1
transform 1 0 22632 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2022
timestamp 1
transform 1 0 27784 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2023
timestamp 1
transform 1 0 32936 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2024
timestamp 1
transform 1 0 38088 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2025
timestamp 1
transform 1 0 43240 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2026
timestamp 1
transform 1 0 48392 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2027
timestamp 1
transform 1 0 53544 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2028
timestamp 1
transform 1 0 58696 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2029
timestamp 1
transform 1 0 63848 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2030
timestamp 1
transform 1 0 69000 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_2031
timestamp 1
transform 1 0 74152 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2032
timestamp 1
transform 1 0 4600 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2033
timestamp 1
transform 1 0 9752 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2034
timestamp 1
transform 1 0 14904 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2035
timestamp 1
transform 1 0 20056 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2036
timestamp 1
transform 1 0 25208 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2037
timestamp 1
transform 1 0 30360 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2038
timestamp 1
transform 1 0 35512 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2039
timestamp 1
transform 1 0 40664 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2040
timestamp 1
transform 1 0 45816 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2041
timestamp 1
transform 1 0 50968 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2042
timestamp 1
transform 1 0 56120 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2043
timestamp 1
transform 1 0 61272 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2044
timestamp 1
transform 1 0 66424 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2045
timestamp 1
transform 1 0 71576 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_2046
timestamp 1
transform 1 0 76728 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2047
timestamp 1
transform 1 0 7176 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2048
timestamp 1
transform 1 0 12328 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2049
timestamp 1
transform 1 0 17480 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2050
timestamp 1
transform 1 0 22632 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2051
timestamp 1
transform 1 0 27784 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2052
timestamp 1
transform 1 0 32936 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2053
timestamp 1
transform 1 0 38088 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2054
timestamp 1
transform 1 0 43240 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2055
timestamp 1
transform 1 0 48392 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2056
timestamp 1
transform 1 0 53544 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2057
timestamp 1
transform 1 0 58696 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2058
timestamp 1
transform 1 0 63848 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2059
timestamp 1
transform 1 0 69000 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_2060
timestamp 1
transform 1 0 74152 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2061
timestamp 1
transform 1 0 4600 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2062
timestamp 1
transform 1 0 9752 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2063
timestamp 1
transform 1 0 14904 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2064
timestamp 1
transform 1 0 20056 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2065
timestamp 1
transform 1 0 25208 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2066
timestamp 1
transform 1 0 30360 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2067
timestamp 1
transform 1 0 35512 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2068
timestamp 1
transform 1 0 40664 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2069
timestamp 1
transform 1 0 45816 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2070
timestamp 1
transform 1 0 50968 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2071
timestamp 1
transform 1 0 56120 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2072
timestamp 1
transform 1 0 61272 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2073
timestamp 1
transform 1 0 66424 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2074
timestamp 1
transform 1 0 71576 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_2075
timestamp 1
transform 1 0 76728 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2076
timestamp 1
transform 1 0 7176 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2077
timestamp 1
transform 1 0 12328 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2078
timestamp 1
transform 1 0 17480 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2079
timestamp 1
transform 1 0 22632 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2080
timestamp 1
transform 1 0 27784 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2081
timestamp 1
transform 1 0 32936 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2082
timestamp 1
transform 1 0 38088 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2083
timestamp 1
transform 1 0 43240 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2084
timestamp 1
transform 1 0 48392 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2085
timestamp 1
transform 1 0 53544 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2086
timestamp 1
transform 1 0 58696 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2087
timestamp 1
transform 1 0 63848 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2088
timestamp 1
transform 1 0 69000 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_2089
timestamp 1
transform 1 0 74152 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2090
timestamp 1
transform 1 0 4600 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2091
timestamp 1
transform 1 0 9752 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2092
timestamp 1
transform 1 0 14904 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2093
timestamp 1
transform 1 0 20056 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2094
timestamp 1
transform 1 0 25208 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2095
timestamp 1
transform 1 0 30360 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2096
timestamp 1
transform 1 0 35512 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2097
timestamp 1
transform 1 0 40664 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2098
timestamp 1
transform 1 0 45816 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2099
timestamp 1
transform 1 0 50968 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2100
timestamp 1
transform 1 0 56120 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2101
timestamp 1
transform 1 0 61272 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2102
timestamp 1
transform 1 0 66424 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2103
timestamp 1
transform 1 0 71576 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_2104
timestamp 1
transform 1 0 76728 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2105
timestamp 1
transform 1 0 7176 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2106
timestamp 1
transform 1 0 12328 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2107
timestamp 1
transform 1 0 17480 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2108
timestamp 1
transform 1 0 22632 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2109
timestamp 1
transform 1 0 27784 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2110
timestamp 1
transform 1 0 32936 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2111
timestamp 1
transform 1 0 38088 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2112
timestamp 1
transform 1 0 43240 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2113
timestamp 1
transform 1 0 48392 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2114
timestamp 1
transform 1 0 53544 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2115
timestamp 1
transform 1 0 58696 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2116
timestamp 1
transform 1 0 63848 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2117
timestamp 1
transform 1 0 69000 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_2118
timestamp 1
transform 1 0 74152 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2119
timestamp 1
transform 1 0 4600 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2120
timestamp 1
transform 1 0 9752 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2121
timestamp 1
transform 1 0 14904 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2122
timestamp 1
transform 1 0 20056 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2123
timestamp 1
transform 1 0 25208 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2124
timestamp 1
transform 1 0 30360 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2125
timestamp 1
transform 1 0 35512 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2126
timestamp 1
transform 1 0 40664 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2127
timestamp 1
transform 1 0 45816 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2128
timestamp 1
transform 1 0 50968 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2129
timestamp 1
transform 1 0 56120 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2130
timestamp 1
transform 1 0 61272 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2131
timestamp 1
transform 1 0 66424 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2132
timestamp 1
transform 1 0 71576 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_2133
timestamp 1
transform 1 0 76728 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2134
timestamp 1
transform 1 0 7176 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2135
timestamp 1
transform 1 0 12328 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2136
timestamp 1
transform 1 0 17480 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2137
timestamp 1
transform 1 0 22632 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2138
timestamp 1
transform 1 0 27784 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2139
timestamp 1
transform 1 0 32936 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2140
timestamp 1
transform 1 0 38088 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2141
timestamp 1
transform 1 0 43240 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2142
timestamp 1
transform 1 0 48392 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2143
timestamp 1
transform 1 0 53544 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2144
timestamp 1
transform 1 0 58696 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2145
timestamp 1
transform 1 0 63848 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2146
timestamp 1
transform 1 0 69000 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_2147
timestamp 1
transform 1 0 74152 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2148
timestamp 1
transform 1 0 4600 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2149
timestamp 1
transform 1 0 9752 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2150
timestamp 1
transform 1 0 14904 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2151
timestamp 1
transform 1 0 20056 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2152
timestamp 1
transform 1 0 25208 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2153
timestamp 1
transform 1 0 30360 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2154
timestamp 1
transform 1 0 35512 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2155
timestamp 1
transform 1 0 40664 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2156
timestamp 1
transform 1 0 45816 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2157
timestamp 1
transform 1 0 50968 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2158
timestamp 1
transform 1 0 56120 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2159
timestamp 1
transform 1 0 61272 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2160
timestamp 1
transform 1 0 66424 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2161
timestamp 1
transform 1 0 71576 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_2162
timestamp 1
transform 1 0 76728 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2163
timestamp 1
transform 1 0 7176 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2164
timestamp 1
transform 1 0 12328 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2165
timestamp 1
transform 1 0 17480 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2166
timestamp 1
transform 1 0 22632 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2167
timestamp 1
transform 1 0 27784 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2168
timestamp 1
transform 1 0 32936 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2169
timestamp 1
transform 1 0 38088 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2170
timestamp 1
transform 1 0 43240 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2171
timestamp 1
transform 1 0 48392 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2172
timestamp 1
transform 1 0 53544 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2173
timestamp 1
transform 1 0 58696 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2174
timestamp 1
transform 1 0 63848 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2175
timestamp 1
transform 1 0 69000 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_2176
timestamp 1
transform 1 0 74152 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2177
timestamp 1
transform 1 0 4600 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2178
timestamp 1
transform 1 0 9752 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2179
timestamp 1
transform 1 0 14904 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2180
timestamp 1
transform 1 0 20056 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2181
timestamp 1
transform 1 0 25208 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2182
timestamp 1
transform 1 0 30360 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2183
timestamp 1
transform 1 0 35512 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2184
timestamp 1
transform 1 0 40664 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2185
timestamp 1
transform 1 0 45816 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2186
timestamp 1
transform 1 0 50968 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2187
timestamp 1
transform 1 0 56120 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2188
timestamp 1
transform 1 0 61272 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2189
timestamp 1
transform 1 0 66424 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2190
timestamp 1
transform 1 0 71576 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_2191
timestamp 1
transform 1 0 76728 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2192
timestamp 1
transform 1 0 7176 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2193
timestamp 1
transform 1 0 12328 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2194
timestamp 1
transform 1 0 17480 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2195
timestamp 1
transform 1 0 22632 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2196
timestamp 1
transform 1 0 27784 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2197
timestamp 1
transform 1 0 32936 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2198
timestamp 1
transform 1 0 38088 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2199
timestamp 1
transform 1 0 43240 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2200
timestamp 1
transform 1 0 48392 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2201
timestamp 1
transform 1 0 53544 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2202
timestamp 1
transform 1 0 58696 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2203
timestamp 1
transform 1 0 63848 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2204
timestamp 1
transform 1 0 69000 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_2205
timestamp 1
transform 1 0 74152 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2206
timestamp 1
transform 1 0 4600 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2207
timestamp 1
transform 1 0 9752 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2208
timestamp 1
transform 1 0 14904 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2209
timestamp 1
transform 1 0 20056 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2210
timestamp 1
transform 1 0 25208 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2211
timestamp 1
transform 1 0 30360 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2212
timestamp 1
transform 1 0 35512 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2213
timestamp 1
transform 1 0 40664 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2214
timestamp 1
transform 1 0 45816 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2215
timestamp 1
transform 1 0 50968 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2216
timestamp 1
transform 1 0 56120 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2217
timestamp 1
transform 1 0 61272 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2218
timestamp 1
transform 1 0 66424 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2219
timestamp 1
transform 1 0 71576 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_2220
timestamp 1
transform 1 0 76728 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2221
timestamp 1
transform 1 0 7176 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2222
timestamp 1
transform 1 0 12328 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2223
timestamp 1
transform 1 0 17480 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2224
timestamp 1
transform 1 0 22632 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2225
timestamp 1
transform 1 0 27784 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2226
timestamp 1
transform 1 0 32936 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2227
timestamp 1
transform 1 0 38088 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2228
timestamp 1
transform 1 0 43240 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2229
timestamp 1
transform 1 0 48392 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2230
timestamp 1
transform 1 0 53544 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2231
timestamp 1
transform 1 0 58696 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2232
timestamp 1
transform 1 0 63848 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2233
timestamp 1
transform 1 0 69000 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_2234
timestamp 1
transform 1 0 74152 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2235
timestamp 1
transform 1 0 4600 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2236
timestamp 1
transform 1 0 9752 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2237
timestamp 1
transform 1 0 14904 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2238
timestamp 1
transform 1 0 20056 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2239
timestamp 1
transform 1 0 25208 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2240
timestamp 1
transform 1 0 30360 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2241
timestamp 1
transform 1 0 35512 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2242
timestamp 1
transform 1 0 40664 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2243
timestamp 1
transform 1 0 45816 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2244
timestamp 1
transform 1 0 50968 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2245
timestamp 1
transform 1 0 56120 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2246
timestamp 1
transform 1 0 61272 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2247
timestamp 1
transform 1 0 66424 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2248
timestamp 1
transform 1 0 71576 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_2249
timestamp 1
transform 1 0 76728 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2250
timestamp 1
transform 1 0 7176 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2251
timestamp 1
transform 1 0 12328 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2252
timestamp 1
transform 1 0 17480 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2253
timestamp 1
transform 1 0 22632 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2254
timestamp 1
transform 1 0 27784 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2255
timestamp 1
transform 1 0 32936 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2256
timestamp 1
transform 1 0 38088 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2257
timestamp 1
transform 1 0 43240 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2258
timestamp 1
transform 1 0 48392 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2259
timestamp 1
transform 1 0 53544 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2260
timestamp 1
transform 1 0 58696 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2261
timestamp 1
transform 1 0 63848 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2262
timestamp 1
transform 1 0 69000 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_2263
timestamp 1
transform 1 0 74152 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2264
timestamp 1
transform 1 0 4600 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2265
timestamp 1
transform 1 0 9752 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2266
timestamp 1
transform 1 0 14904 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2267
timestamp 1
transform 1 0 20056 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2268
timestamp 1
transform 1 0 25208 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2269
timestamp 1
transform 1 0 30360 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2270
timestamp 1
transform 1 0 35512 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2271
timestamp 1
transform 1 0 40664 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2272
timestamp 1
transform 1 0 45816 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2273
timestamp 1
transform 1 0 50968 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2274
timestamp 1
transform 1 0 56120 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2275
timestamp 1
transform 1 0 61272 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2276
timestamp 1
transform 1 0 66424 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2277
timestamp 1
transform 1 0 71576 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_2278
timestamp 1
transform 1 0 76728 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2279
timestamp 1
transform 1 0 7176 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2280
timestamp 1
transform 1 0 12328 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2281
timestamp 1
transform 1 0 17480 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2282
timestamp 1
transform 1 0 22632 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2283
timestamp 1
transform 1 0 27784 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2284
timestamp 1
transform 1 0 32936 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2285
timestamp 1
transform 1 0 38088 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2286
timestamp 1
transform 1 0 43240 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2287
timestamp 1
transform 1 0 48392 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2288
timestamp 1
transform 1 0 53544 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2289
timestamp 1
transform 1 0 58696 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2290
timestamp 1
transform 1 0 63848 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2291
timestamp 1
transform 1 0 69000 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_2292
timestamp 1
transform 1 0 74152 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2293
timestamp 1
transform 1 0 4600 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2294
timestamp 1
transform 1 0 7176 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2295
timestamp 1
transform 1 0 9752 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2296
timestamp 1
transform 1 0 12328 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2297
timestamp 1
transform 1 0 14904 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2298
timestamp 1
transform 1 0 17480 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2299
timestamp 1
transform 1 0 20056 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2300
timestamp 1
transform 1 0 22632 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2301
timestamp 1
transform 1 0 25208 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2302
timestamp 1
transform 1 0 27784 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2303
timestamp 1
transform 1 0 30360 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2304
timestamp 1
transform 1 0 32936 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2305
timestamp 1
transform 1 0 35512 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2306
timestamp 1
transform 1 0 38088 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2307
timestamp 1
transform 1 0 40664 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2308
timestamp 1
transform 1 0 43240 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2309
timestamp 1
transform 1 0 45816 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2310
timestamp 1
transform 1 0 48392 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2311
timestamp 1
transform 1 0 50968 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2312
timestamp 1
transform 1 0 53544 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2313
timestamp 1
transform 1 0 56120 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2314
timestamp 1
transform 1 0 58696 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2315
timestamp 1
transform 1 0 61272 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2316
timestamp 1
transform 1 0 63848 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2317
timestamp 1
transform 1 0 66424 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2318
timestamp 1
transform 1 0 69000 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2319
timestamp 1
transform 1 0 71576 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2320
timestamp 1
transform 1 0 74152 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_2321
timestamp 1
transform 1 0 76728 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  TopModule_7
timestamp 1
transform -1 0 2576 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_8
timestamp 1
transform -1 0 49956 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_9
timestamp 1
transform 1 0 77372 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_10
timestamp 1
transform -1 0 33304 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_11
timestamp 1
transform -1 0 59616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_12
timestamp 1
transform 1 0 77372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_13
timestamp 1
transform -1 0 2576 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_14
timestamp 1
transform -1 0 42228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_15
timestamp 1
transform -1 0 59064 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_16
timestamp 1
transform -1 0 2576 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_17
timestamp 1
transform -1 0 2576 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_18
timestamp 1
transform -1 0 52532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_19
timestamp 1
transform -1 0 2576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_20
timestamp 1
transform -1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_21
timestamp 1
transform 1 0 77372 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_22
timestamp 1
transform -1 0 58328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_23
timestamp 1
transform -1 0 2576 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_24
timestamp 1
transform -1 0 24196 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_25
timestamp 1
transform -1 0 2576 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_26
timestamp 1
transform -1 0 2576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_27
timestamp 1
transform -1 0 40296 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_28
timestamp 1
transform -1 0 54464 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_29
timestamp 1
transform -1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_30
timestamp 1
transform 1 0 77372 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_31
timestamp 1
transform -1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_32
timestamp 1
transform -1 0 44804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_33
timestamp 1
transform -1 0 42872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  TopModule_34
timestamp 1
transform -1 0 42228 0 1 77248
box -38 -48 314 592
<< labels >>
flabel metal4 s 5788 2128 6108 77840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 36508 2128 36828 77840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 67228 2128 67548 77840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1976 6006 77972 6326 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1976 36642 77972 36962 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1976 67278 77972 67598 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5128 2128 5448 77840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 35848 2128 36168 77840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 66568 2128 66888 77840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1976 5346 77972 5666 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1976 35982 77972 36302 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1976 66618 77972 66938 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 ctrl[0]
port 3 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 ctrl[1]
port 4 nsew signal input
flabel metal3 s 79200 38768 80000 38888 0 FreeSans 480 0 0 0 data_out[0]
port 5 nsew signal output
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 data_out[10]
port 6 nsew signal output
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 data_out[11]
port 7 nsew signal output
flabel metal2 s 58622 79200 58678 80000 0 FreeSans 224 90 0 0 data_out[12]
port 8 nsew signal output
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 data_out[13]
port 9 nsew signal output
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 data_out[14]
port 10 nsew signal output
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 data_out[15]
port 11 nsew signal output
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 data_out[16]
port 12 nsew signal output
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 data_out[17]
port 13 nsew signal output
flabel metal3 s 79200 51688 80000 51808 0 FreeSans 480 0 0 0 data_out[18]
port 14 nsew signal output
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 data_out[19]
port 15 nsew signal output
flabel metal3 s 79200 37408 80000 37528 0 FreeSans 480 0 0 0 data_out[1]
port 16 nsew signal output
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 data_out[20]
port 17 nsew signal output
flabel metal2 s 23846 79200 23902 80000 0 FreeSans 224 90 0 0 data_out[21]
port 18 nsew signal output
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 data_out[22]
port 19 nsew signal output
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 data_out[23]
port 20 nsew signal output
flabel metal2 s 39946 79200 40002 80000 0 FreeSans 224 90 0 0 data_out[24]
port 21 nsew signal output
flabel metal2 s 54114 79200 54170 80000 0 FreeSans 224 90 0 0 data_out[25]
port 22 nsew signal output
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 data_out[26]
port 23 nsew signal output
flabel metal3 s 79200 21088 80000 21208 0 FreeSans 480 0 0 0 data_out[27]
port 24 nsew signal output
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 data_out[28]
port 25 nsew signal output
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 data_out[29]
port 26 nsew signal output
flabel metal3 s 79200 36728 80000 36848 0 FreeSans 480 0 0 0 data_out[2]
port 27 nsew signal output
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 data_out[30]
port 28 nsew signal output
flabel metal2 s 41878 79200 41934 80000 0 FreeSans 224 90 0 0 data_out[31]
port 29 nsew signal output
flabel metal3 s 79200 38088 80000 38208 0 FreeSans 480 0 0 0 data_out[3]
port 30 nsew signal output
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 data_out[4]
port 31 nsew signal output
flabel metal2 s 49606 79200 49662 80000 0 FreeSans 224 90 0 0 data_out[5]
port 32 nsew signal output
flabel metal3 s 79200 49648 80000 49768 0 FreeSans 480 0 0 0 data_out[6]
port 33 nsew signal output
flabel metal2 s 32862 79200 32918 80000 0 FreeSans 224 90 0 0 data_out[7]
port 34 nsew signal output
flabel metal2 s 59266 0 59322 800 0 FreeSans 224 90 0 0 data_out[8]
port 35 nsew signal output
flabel metal3 s 79200 16328 80000 16448 0 FreeSans 480 0 0 0 data_out[9]
port 36 nsew signal output
flabel metal3 s 79200 34008 80000 34128 0 FreeSans 480 0 0 0 reset
port 37 nsew signal input
rlabel metal1 39974 77248 39974 77248 0 VGND
rlabel metal1 39974 77792 39974 77792 0 VPWR
rlabel metal2 58926 42466 58926 42466 0 _000_
rlabel metal1 58519 39338 58519 39338 0 _001_
rlabel metal1 58059 34986 58059 34986 0 _002_
rlabel metal1 62107 35734 62107 35734 0 _003_
rlabel metal1 62008 40018 62008 40018 0 _004_
rlabel metal1 66891 43350 66891 43350 0 _005_
rlabel metal1 67114 40018 67114 40018 0 _006_
rlabel metal1 66056 36890 66056 36890 0 _007_
rlabel metal2 66930 33796 66930 33796 0 _008_
rlabel metal1 70656 34170 70656 34170 0 _009_
rlabel metal1 75861 36074 75861 36074 0 _010_
rlabel metal2 71254 41310 71254 41310 0 _011_
rlabel metal1 76091 41514 76091 41514 0 _012_
rlabel metal1 75394 38522 75394 38522 0 _013_
rlabel metal1 75670 38726 75670 38726 0 _014_
rlabel metal2 71622 39202 71622 39202 0 _015_
rlabel metal1 57224 37094 57224 37094 0 _016_
rlabel metal1 57270 38284 57270 38284 0 _017_
rlabel metal2 64630 40868 64630 40868 0 _018_
rlabel metal1 60582 36278 60582 36278 0 _019_
rlabel metal2 64906 42806 64906 42806 0 _020_
rlabel metal1 65734 39814 65734 39814 0 _021_
rlabel metal1 66516 39882 66516 39882 0 _022_
rlabel metal1 66930 36142 66930 36142 0 _023_
rlabel metal1 66148 36346 66148 36346 0 _024_
rlabel metal1 71668 35598 71668 35598 0 _025_
rlabel metal1 70978 38930 70978 38930 0 _026_
rlabel metal1 72220 36210 72220 36210 0 _027_
rlabel metal2 71162 40800 71162 40800 0 _028_
rlabel metal2 71530 39848 71530 39848 0 _029_
rlabel metal1 75578 38862 75578 38862 0 aluop\[0\]
rlabel metal2 74658 38624 74658 38624 0 aluop\[1\]
rlabel metal2 75946 40052 75946 40052 0 aluop\[2\]
rlabel metal3 1004 45628 1004 45628 0 clk
rlabel metal1 66608 38726 66608 38726 0 clknet_0_clk
rlabel metal1 57224 39474 57224 39474 0 clknet_1_0__leaf_clk
rlabel metal1 70242 41174 70242 41174 0 clknet_1_1__leaf_clk
rlabel via2 77510 38811 77510 38811 0 data_out[0]
rlabel metal2 77510 37553 77510 37553 0 data_out[1]
rlabel metal2 77510 36941 77510 36941 0 data_out[2]
rlabel via2 77510 38165 77510 38165 0 data_out[3]
rlabel metal2 70702 35292 70702 35292 0 instruction\[10\]
rlabel metal2 70150 35054 70150 35054 0 instruction\[11\]
rlabel metal1 59754 42738 59754 42738 0 instruction\[2\]
rlabel metal2 60214 36482 60214 36482 0 instruction\[3\]
rlabel metal2 60306 36482 60306 36482 0 instruction\[4\]
rlabel metal1 60030 36108 60030 36108 0 instruction\[5\]
rlabel metal2 64814 41038 64814 41038 0 instruction\[6\]
rlabel metal2 66930 43588 66930 43588 0 instruction\[7\]
rlabel metal1 66746 40630 66746 40630 0 instruction\[8\]
rlabel metal1 67022 37230 67022 37230 0 instruction\[9\]
rlabel metal1 76406 41616 76406 41616 0 net1
rlabel metal1 32982 77690 32982 77690 0 net10
rlabel metal2 59294 1588 59294 1588 0 net11
rlabel metal3 78484 16388 78484 16388 0 net12
rlabel metal3 1510 25908 1510 25908 0 net13
rlabel metal2 41906 1588 41906 1588 0 net14
rlabel metal1 58742 77690 58742 77690 0 net15
rlabel metal3 958 32028 958 32028 0 net16
rlabel metal3 958 27948 958 27948 0 net17
rlabel metal2 52210 1588 52210 1588 0 net18
rlabel metal3 1510 23188 1510 23188 0 net19
rlabel metal2 76314 38726 76314 38726 0 net2
rlabel metal2 33534 1588 33534 1588 0 net20
rlabel via2 77602 51765 77602 51765 0 net21
rlabel metal2 58006 1588 58006 1588 0 net22
rlabel metal3 958 35428 958 35428 0 net23
rlabel metal1 23920 77690 23920 77690 0 net24
rlabel metal3 958 41548 958 41548 0 net25
rlabel metal3 958 26588 958 26588 0 net26
rlabel metal1 40020 77690 40020 77690 0 net27
rlabel metal1 54188 77690 54188 77690 0 net28
rlabel metal2 23230 1588 23230 1588 0 net29
rlabel metal2 76498 37094 76498 37094 0 net3
rlabel metal2 77602 21233 77602 21233 0 net30
rlabel metal2 22586 1588 22586 1588 0 net31
rlabel metal2 44482 1588 44482 1588 0 net32
rlabel metal2 42550 1588 42550 1588 0 net33
rlabel metal1 41952 77690 41952 77690 0 net34
rlabel metal1 58190 42228 58190 42228 0 net35
rlabel metal1 74888 41106 74888 41106 0 net36
rlabel metal1 65918 36788 65918 36788 0 net37
rlabel metal1 57086 35666 57086 35666 0 net38
rlabel metal1 66148 34578 66148 34578 0 net39
rlabel metal1 76314 37162 76314 37162 0 net4
rlabel metal1 65780 43758 65780 43758 0 net40
rlabel metal1 73002 36142 73002 36142 0 net41
rlabel metal1 61456 40154 61456 40154 0 net42
rlabel metal1 70886 35598 70886 35598 0 net43
rlabel metal1 76820 38318 76820 38318 0 net5
rlabel metal1 58604 39406 58604 39406 0 net6
rlabel metal3 1510 28628 1510 28628 0 net7
rlabel metal1 49680 77690 49680 77690 0 net8
rlabel via2 77602 49725 77602 49725 0 net9
rlabel metal2 77510 34323 77510 34323 0 reset
rlabel metal2 68034 34204 68034 34204 0 u_pc.next_pc\[10\]
rlabel metal2 71346 35054 71346 35054 0 u_pc.next_pc\[11\]
rlabel metal1 74382 36040 74382 36040 0 u_pc.next_pc\[12\]
rlabel metal1 70610 40698 70610 40698 0 u_pc.next_pc\[13\]
rlabel metal1 74750 41038 74750 41038 0 u_pc.next_pc\[14\]
rlabel metal1 58052 42330 58052 42330 0 u_pc.next_pc\[2\]
rlabel metal2 57086 38930 57086 38930 0 u_pc.next_pc\[3\]
rlabel metal1 56524 35258 56524 35258 0 u_pc.next_pc\[4\]
rlabel metal1 60628 35734 60628 35734 0 u_pc.next_pc\[5\]
rlabel metal1 61446 40698 61446 40698 0 u_pc.next_pc\[6\]
rlabel metal2 65458 43486 65458 43486 0 u_pc.next_pc\[7\]
rlabel metal1 67390 40154 67390 40154 0 u_pc.next_pc\[8\]
rlabel metal1 65412 36890 65412 36890 0 u_pc.next_pc\[9\]
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>
