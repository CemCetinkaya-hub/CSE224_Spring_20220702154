* NGSPICE file created from TopModule.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

.subckt TopModule VGND VPWR clk ctrl[0] ctrl[1] data_out[0] data_out[10] data_out[11]
+ data_out[12] data_out[13] data_out[14] data_out[15] data_out[16] data_out[17] data_out[18]
+ data_out[19] data_out[1] data_out[20] data_out[21] data_out[22] data_out[23] data_out[24]
+ data_out[25] data_out[26] data_out[27] data_out[28] data_out[29] data_out[2] data_out[30]
+ data_out[31] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7] data_out[8]
+ data_out[9] reset
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_062_ net36 _028_ VGND VGND VPWR VPWR u_pc.next_pc\[14\] sky130_fd_sc_hd__xor2_1
XFILLER_137_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_045_ net42 _018_ VGND VGND VPWR VPWR u_pc.next_pc\[6\] sky130_fd_sc_hd__xor2_1
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_061_ _028_ _029_ VGND VGND VPWR VPWR u_pc.next_pc\[13\] sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_044_ instruction\[6\] _018_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__nand2_1
XFILLER_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_060_ aluop\[0\] _018_ _023_ _026_ aluop\[1\] VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__a41o_1
XFILLER_136_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_043_ _018_ _019_ VGND VGND VPWR VPWR u_pc.next_pc\[5\] sky130_fd_sc_hd__and2b_1
XFILLER_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_121_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_042_ instruction\[2\] instruction\[3\] instruction\[4\] instruction\[5\] VGND VGND
+ VPWR VPWR _019_ sky130_fd_sc_hd__a31o_1
XFILLER_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 clknet_1_1__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_041_ instruction\[2\] instruction\[3\] instruction\[4\] instruction\[5\] VGND VGND
+ VPWR VPWR _018_ sky130_fd_sc_hd__and4_4
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_26_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_040_ net38 _016_ VGND VGND VPWR VPWR u_pc.next_pc\[4\] sky130_fd_sc_hd__xnor2_1
XFILLER_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_119_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_15_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_31_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_86_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_95_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_079_ clknet_1_0__leaf_clk u_pc.next_pc\[6\] _004_ VGND VGND VPWR VPWR instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_124_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_078_ clknet_1_0__leaf_clk u_pc.next_pc\[5\] _003_ VGND VGND VPWR VPWR instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_112_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_077_ clknet_1_0__leaf_clk u_pc.next_pc\[4\] _002_ VGND VGND VPWR VPWR instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_29_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_56_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_91_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 reset VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_84_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_7 VGND VGND VPWR VPWR TopModule_7/HI data_out[4] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_69_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_076_ clknet_1_0__leaf_clk u_pc.next_pc\[3\] _001_ VGND VGND VPWR VPWR instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_124_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_102_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_059_ _015_ _018_ _023_ _026_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_55_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_8 VGND VGND VPWR VPWR TopModule_8/HI data_out[5] sky130_fd_sc_hd__conb_1
XFILLER_36_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_075_ clknet_1_0__leaf_clk u_pc.next_pc\[2\] _000_ VGND VGND VPWR VPWR instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_124_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_058_ net41 _027_ VGND VGND VPWR VPWR u_pc.next_pc\[12\] sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_55_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_9 VGND VGND VPWR VPWR TopModule_9/HI data_out[6] sky130_fd_sc_hd__conb_1
XFILLER_36_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_074_ net1 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__inv_2
XFILLER_109_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_25_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_057_ _025_ _027_ VGND VGND VPWR VPWR u_pc.next_pc\[11\] sky130_fd_sc_hd__and2_1
XFILLER_124_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_073_ net1 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__inv_2
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_056_ _018_ _023_ _026_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__nand3_1
XFILLER_124_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_039_ _016_ _017_ VGND VGND VPWR VPWR u_pc.next_pc\[3\] sky130_fd_sc_hd__and2_1
XFILLER_125_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_118_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_072_ net1 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
XFILLER_137_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_055_ instruction\[10\] instruction\[11\] VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and2_1
XFILLER_124_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_038_ instruction\[2\] instruction\[3\] VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__or2_1
XFILLER_125_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_071_ net6 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__inv_2
XFILLER_136_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_054_ instruction\[10\] _018_ _023_ net43 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_12_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_037_ instruction\[2\] instruction\[3\] VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__nand2_1
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_070_ net6 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__inv_2
XFILLER_136_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_053_ net39 _024_ VGND VGND VPWR VPWR u_pc.next_pc\[10\] sky130_fd_sc_hd__xnor2_1
XFILLER_137_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_036_ _013_ aluop\[0\] _014_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__a21oi_1
XFILLER_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_123_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_052_ net37 _021_ _024_ VGND VGND VPWR VPWR u_pc.next_pc\[9\] sky130_fd_sc_hd__o21a_1
XFILLER_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_035_ aluop\[1\] aluop\[0\] VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__and2_1
XFILLER_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_051_ _018_ _023_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__nand2_1
XFILLER_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_034_ _014_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__inv_2
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1 instruction\[2\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_683 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_050_ instruction\[6\] instruction\[7\] instruction\[8\] instruction\[9\] VGND VGND
+ VPWR VPWR _023_ sky130_fd_sc_hd__and4_1
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_033_ aluop\[1\] aluop\[2\] aluop\[0\] VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__mux2_1
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2 aluop\[2\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_101_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_032_ net6 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__inv_2
XFILLER_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3 instruction\[9\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_728 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_031_ net35 VGND VGND VPWR VPWR u_pc.next_pc\[2\] sky130_fd_sc_hd__inv_2
XFILLER_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 instruction\[4\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_30 VGND VGND VPWR VPWR TopModule_30/HI data_out[27] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_108_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_030_ aluop\[1\] VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__inv_2
XFILLER_20_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 instruction\[10\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_79_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_97_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTopModule_20 VGND VGND VPWR VPWR TopModule_20/HI data_out[17] sky130_fd_sc_hd__conb_1
XTopModule_31 VGND VGND VPWR VPWR TopModule_31/HI data_out[28] sky130_fd_sc_hd__conb_1
XFILLER_55_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_117_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_126_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 instruction\[7\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_59_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_10 VGND VGND VPWR VPWR TopModule_10/HI data_out[7] sky130_fd_sc_hd__conb_1
XTopModule_21 VGND VGND VPWR VPWR TopModule_21/HI data_out[18] sky130_fd_sc_hd__conb_1
XFILLER_55_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_32 VGND VGND VPWR VPWR TopModule_32/HI data_out[29] sky130_fd_sc_hd__conb_1
XFILLER_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold7 aluop\[0\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTopModule_22 VGND VGND VPWR VPWR TopModule_22/HI data_out[19] sky130_fd_sc_hd__conb_1
XTopModule_11 VGND VGND VPWR VPWR TopModule_11/HI data_out[8] sky130_fd_sc_hd__conb_1
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_33 VGND VGND VPWR VPWR TopModule_33/HI data_out[30] sky130_fd_sc_hd__conb_1
XFILLER_63_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_087_ clknet_1_1__leaf_clk u_pc.next_pc\[14\] _012_ VGND VGND VPWR VPWR aluop\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 instruction\[6\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_128_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_12 VGND VGND VPWR VPWR TopModule_12/HI data_out[9] sky130_fd_sc_hd__conb_1
XTopModule_34 VGND VGND VPWR VPWR TopModule_34/HI data_out[31] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_108_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTopModule_23 VGND VGND VPWR VPWR TopModule_23/HI data_out[20] sky130_fd_sc_hd__conb_1
XFILLER_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_086_ clknet_1_1__leaf_clk u_pc.next_pc\[13\] _011_ VGND VGND VPWR VPWR aluop\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_104_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 instruction\[11\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_113_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_122_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_069_ net6 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__inv_2
XFILLER_112_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_13 VGND VGND VPWR VPWR TopModule_13/HI data_out[10] sky130_fd_sc_hd__conb_1
XFILLER_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTopModule_24 VGND VGND VPWR VPWR TopModule_24/HI data_out[21] sky130_fd_sc_hd__conb_1
XFILLER_64_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_085_ clknet_1_1__leaf_clk u_pc.next_pc\[12\] _010_ VGND VGND VPWR VPWR aluop\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_124_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_068_ net6 VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__inv_2
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTopModule_25 VGND VGND VPWR VPWR TopModule_25/HI data_out[22] sky130_fd_sc_hd__conb_1
XFILLER_64_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_14 VGND VGND VPWR VPWR TopModule_14/HI data_out[11] sky130_fd_sc_hd__conb_1
XFILLER_36_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_084_ clknet_1_1__leaf_clk u_pc.next_pc\[11\] _009_ VGND VGND VPWR VPWR instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_067_ net6 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__inv_2
XFILLER_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput2 net2 VGND VGND VPWR VPWR data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_15 VGND VGND VPWR VPWR TopModule_15/HI data_out[12] sky130_fd_sc_hd__conb_1
XFILLER_64_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTopModule_26 VGND VGND VPWR VPWR TopModule_26/HI data_out[23] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_108_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_083_ clknet_1_1__leaf_clk u_pc.next_pc\[10\] _008_ VGND VGND VPWR VPWR instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_124_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_066_ net6 VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__inv_2
XFILLER_124_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_049_ _021_ _022_ VGND VGND VPWR VPWR u_pc.next_pc\[8\] sky130_fd_sc_hd__and2b_1
XFILLER_125_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput3 net3 VGND VGND VPWR VPWR data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_110_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_27 VGND VGND VPWR VPWR TopModule_27/HI data_out[24] sky130_fd_sc_hd__conb_1
XFILLER_64_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_16 VGND VGND VPWR VPWR TopModule_16/HI data_out[13] sky130_fd_sc_hd__conb_1
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_90_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_082_ clknet_1_0__leaf_clk u_pc.next_pc\[9\] _007_ VGND VGND VPWR VPWR instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_065_ net6 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__inv_2
XFILLER_124_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_117_ net5 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_048_ instruction\[6\] instruction\[7\] _018_ instruction\[8\] VGND VGND VPWR VPWR
+ _022_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_59_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_110_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_721 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput4 net4 VGND VGND VPWR VPWR data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_96_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_28 VGND VGND VPWR VPWR TopModule_28/HI data_out[25] sky130_fd_sc_hd__conb_1
XTopModule_17 VGND VGND VPWR VPWR TopModule_17/HI data_out[14] sky130_fd_sc_hd__conb_1
XFILLER_64_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_113_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_081_ clknet_1_1__leaf_clk u_pc.next_pc\[8\] _006_ VGND VGND VPWR VPWR instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_064_ net6 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__inv_2
XFILLER_124_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_116_ net4 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_047_ instruction\[6\] instruction\[7\] instruction\[8\] _018_ VGND VGND VPWR VPWR
+ _021_ sky130_fd_sc_hd__and4_1
XFILLER_124_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput5 net5 VGND VGND VPWR VPWR data_out[3] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTopModule_29 VGND VGND VPWR VPWR TopModule_29/HI data_out[26] sky130_fd_sc_hd__conb_1
XTopModule_18 VGND VGND VPWR VPWR TopModule_18/HI data_out[15] sky130_fd_sc_hd__conb_1
XFILLER_48_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_080_ clknet_1_0__leaf_clk u_pc.next_pc\[7\] _005_ VGND VGND VPWR VPWR instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_87_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_063_ net6 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
XFILLER_137_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_046_ net40 _020_ VGND VGND VPWR VPWR u_pc.next_pc\[7\] sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_59_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout6 net1 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTopModule_19 VGND VGND VPWR VPWR TopModule_19/HI data_out[16] sky130_fd_sc_hd__conb_1
XFILLER_48_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

